magic
tech scmos
timestamp 1731058680
<< nwell >>
rect -186 0 -162 56
rect -153 0 -129 56
rect -120 0 -96 56
rect -87 0 -63 56
rect -54 0 -30 56
rect -16 0 8 56
<< polysilicon >>
rect -175 50 -173 53
rect -142 50 -140 53
rect -109 50 -107 53
rect -76 50 -74 53
rect -43 50 -41 53
rect -5 50 -3 53
rect -175 -3 -173 10
rect -142 -3 -140 10
rect -109 -3 -107 10
rect -76 -3 -74 10
rect -43 -3 -41 10
rect -5 -12 -3 10
rect -67 -33 -64 -31
rect -24 -33 -21 -31
rect -5 -35 -3 -32
rect -67 -52 -64 -50
rect -24 -52 -21 -50
rect -67 -71 -64 -69
rect -24 -71 -21 -69
rect -67 -90 -64 -88
rect -24 -90 -21 -88
rect -67 -109 -64 -107
rect -24 -109 -21 -107
<< ndiffusion >>
rect -64 -31 -24 -30
rect -6 -32 -5 -12
rect -3 -32 -2 -12
rect -64 -34 -24 -33
rect -64 -50 -24 -49
rect -64 -53 -24 -52
rect -64 -69 -24 -68
rect -64 -72 -24 -71
rect -64 -88 -24 -87
rect -64 -91 -24 -90
rect -64 -107 -24 -106
rect -64 -110 -24 -109
<< pdiffusion >>
rect -176 10 -175 50
rect -173 10 -172 50
rect -143 10 -142 50
rect -140 10 -139 50
rect -110 10 -109 50
rect -107 10 -106 50
rect -77 10 -76 50
rect -74 10 -73 50
rect -44 10 -43 50
rect -41 10 -40 50
rect -6 10 -5 50
rect -3 10 -2 50
<< metal1 >>
rect -186 60 8 63
rect -186 56 -162 60
rect -153 56 -129 60
rect -120 56 -96 60
rect -87 56 -63 60
rect -54 56 -30 60
rect -16 56 8 60
rect -180 50 -176 56
rect -147 50 -143 56
rect -114 50 -110 56
rect -81 50 -77 56
rect -48 50 -44 56
rect -10 50 -6 56
rect -172 0 -168 10
rect -139 0 -135 10
rect -106 0 -102 10
rect -73 0 -69 10
rect -40 0 -36 10
rect -176 -105 -172 -7
rect -143 -86 -139 -7
rect -110 -67 -106 -7
rect -87 -7 -77 -3
rect -2 -4 2 10
rect -87 -48 -83 -7
rect -44 -12 -40 -7
rect -73 -15 -40 -12
rect -28 -8 -9 -4
rect -2 -8 13 -4
rect -73 -29 -67 -15
rect -28 -26 -24 -8
rect -2 -12 2 -8
rect -10 -34 -6 -32
rect -28 -45 -24 -38
rect -87 -54 -73 -48
rect -16 -37 -6 -34
rect -28 -64 -24 -57
rect -110 -73 -73 -67
rect -28 -83 -24 -76
rect -143 -92 -73 -86
rect -28 -102 -24 -95
rect -176 -111 -73 -105
rect -16 -110 -12 -37
rect -24 -114 -12 -110
<< metal2 >>
rect -168 0 -139 5
rect -135 0 -106 5
rect -102 0 -73 5
rect -69 0 -40 5
rect -36 0 -19 5
rect -23 -4 -19 0
<< ntransistor >>
rect -64 -33 -24 -31
rect -5 -32 -3 -12
rect -64 -52 -24 -50
rect -64 -71 -24 -69
rect -64 -90 -24 -88
rect -64 -109 -24 -107
<< ptransistor >>
rect -175 10 -173 50
rect -142 10 -140 50
rect -109 10 -107 50
rect -76 10 -74 50
rect -43 10 -41 50
rect -5 10 -3 50
<< polycontact >>
rect -176 -7 -172 -3
rect -143 -7 -139 -3
rect -110 -7 -106 -3
rect -77 -7 -73 -3
rect -44 -7 -40 -3
rect -9 -8 -5 -4
rect -73 -35 -67 -29
rect -73 -54 -67 -48
rect -73 -73 -67 -67
rect -73 -92 -67 -86
rect -73 -111 -67 -105
<< ndcontact >>
rect -64 -30 -24 -26
rect -10 -32 -6 -12
rect -2 -32 2 -12
rect -64 -38 -24 -34
rect -64 -49 -24 -45
rect -64 -57 -24 -53
rect -64 -68 -24 -64
rect -64 -76 -24 -72
rect -64 -87 -24 -83
rect -64 -95 -24 -91
rect -64 -106 -24 -102
rect -64 -114 -24 -110
<< pdcontact >>
rect -180 10 -176 50
rect -172 10 -168 50
rect -147 10 -143 50
rect -139 10 -135 50
rect -114 10 -110 50
rect -106 10 -102 50
rect -81 10 -77 50
rect -73 10 -69 50
rect -48 10 -44 50
rect -40 10 -36 50
rect -10 10 -6 50
rect -2 10 2 50
<< pad >>
rect -172 0 -168 5
rect -139 0 -135 5
rect -106 0 -102 5
rect -73 0 -69 5
rect -40 0 -36 5
rect -23 -8 -19 -4
<< labels >>
rlabel metal1 -15 -6 -15 -6 1 ybar
rlabel metal1 -109 -11 -109 -11 1 a
rlabel metal1 -42 -12 -42 -12 1 c
rlabel metal1 -53 62 -53 62 5 vdd
rlabel metal1 -82 -5 -82 -5 1 b
rlabel metal1 -15 -74 -15 -74 1 gnd
rlabel metal1 6 -6 6 -6 1 y
rlabel metal1 -142 -12 -142 -12 1 d
rlabel metal1 -174 -12 -174 -12 1 e
<< end >>
