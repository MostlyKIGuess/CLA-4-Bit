magic
tech scmos
timestamp 1731868666
use testing  testing_0
timestamp 1731837759
transform 1 0 129 0 1 474
box -129 -474 1258 717
<< end >>
