* SPICE3 file created from cla.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Power Supply for the circuit
Vdd vdd gnd 'SUPPLY'


* Input Signals
* for testing
* Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
* Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 30n 60n)     
* Va1 a1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 10n 20n)    
* Vb1 b1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 30n 60n)    
* Va2 a2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 10n 20n)   
* Vb2 b2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 30n 60n)   
* Va3 a3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 10n 20n)   
* Vb3 b3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 30n 60n)   
* Vcin cin gnd DC 0         

* Input Signals for delay measurement

*  falling and rising
Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
Va1 a1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
Vb1 b1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
Va2 a2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Vb2 b2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Va3 a3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Vb3 b3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Vcin cin gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)

* SPICE3 file created from testing.ext - technology: scmos

.option scale=90n

M1000 a_594_537# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1001 a_239_604# p3 g2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_329_n305# a_325_n314# p3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 a_218_418# p2 vdd w_205_450# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_825_350# g3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 a_600_239# p1p0c0 a_617_278# w_611_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 s1 p1 c1 w_818_n75# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 c1 a_445_147# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1008 p3p2p1g0 a_518_635# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1009 a_693_378# p2g1 a_731_417# w_725_411# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_564_n251# a2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1011 a_600_239# p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 a_594_n65# a1 b1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 gnd a_269_20# p0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 a_594_556# p2 a_594_537# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 a_445_147# g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1016 a_594_575# p1 a_594_556# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1017 p2g1 a_327_429# vdd w_347_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1018 a_440_412# p1 a_440_393# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_564_n389# a3 vdd w_551_n357# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1020 p1p0c0 a_453_311# vdd w_544_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1021 a3 b3 p3 w_329_n384# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 a_518_635# p3 vdd w_505_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a_731_457# p2p1p0c0 a_731_417# w_725_444# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1024 a_808_n381# p3 vdd w_795_n349# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1025 b2 a2 p2 w_368_n246# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1026 p3p2g1 a_381_614# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 p2p1p0c0 a_534_474# vdd w_658_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1028 a_610_395# p1 a_610_377# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1029 a_329_n171# a_325_n180# p2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 a_518_635# g0 a_594_575# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 s2 a_795_n247# a_873_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 vdd a0 a_324_88# w_400_28# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1033 a_594_n65# a_561_n113# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1034 vdd a_302_20# a_269_20# w_291_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 a_325_n180# b2 p2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 a_825_350# p3p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1037 a_304_190# a_271_142# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1038 a_847_245# a_771_282# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1039 a_884_498# p3g2 a_883_464# w_878_485# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 a_731_492# p2p1g0 a_731_457# w_725_479# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1041 a_673_n378# a_597_n341# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 a_597_n341# a_564_n389# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1043 a_315_567# a_239_604# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 g0 a_673_36# vdd w_693_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 p3g2 a_315_567# vdd w_335_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 vdd g3 a_884_498# w_879_518# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1047 a_825_350# p3p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 pocin a_380_153# vdd w_400_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 vdd a_269_20# p0 w_258_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 a_218_418# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1051 a_380_153# a_304_190# vdd w_367_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 b1 a1 a_302_n114# w_367_n112# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_825_350# p3p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1054 a_271_280# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1055 p3p2p1g0 a_518_635# vdd w_642_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_239_604# a_206_556# g2 w_226_594# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 a_304_190# a_271_142# cin w_291_180# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 c3 a_693_378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 g3 a_673_n378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 p2p1g0 a_397_472# vdd w_488_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_440_393# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_688_664# p0 vdd w_774_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 s2 p2 c2 w_815_n209# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1064 a_445_147# pocin gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 p2g1 a_327_429# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 a_600_239# p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1067 a_795_n247# p2 vdd w_782_n215# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_564_n251# a2 vdd w_551_n219# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_327_429# a_251_466# vdd w_314_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 a_688_664# cin vdd w_807_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1071 a_693_378# p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_251_466# p2 g1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 s1 c1 a_798_n113# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_798_n113# p1 vdd w_785_n81# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_325_n314# b3 p3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 a_738_234# p0 vdd w_725_266# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1077 a_673_36# a_597_73# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1078 a_564_25# a0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1079 p3p2g1 a_381_614# vdd w_472_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1080 a_597_n341# a_564_n389# b3 w_584_n351# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1081 a_206_556# p3 vdd w_193_588# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_424_535# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1083 g2 a_564_n251# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1084 g1 a_670_n102# vdd w_690_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1085 s3 p3 c3 w_828_n343# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_610_377# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1087 s0 a_847_245# vdd w_867_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1088 vdd a2 a_325_n180# w_401_n240# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_670_n102# a_594_n65# vdd w_657_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 c4 a_825_350# vdd w_942_382# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_670_n102# a_594_n65# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_424_554# p2 a_424_535# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 a_453_311# p0 vdd w_473_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1094 a_315_567# a_239_604# vdd w_302_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 p3p2p1p0c0 a_688_664# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_771_282# p0 cin w_758_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1097 s1 c1 p1 w_857_n67# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_271_142# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1099 a_534_474# cin vdd w_620_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_534_474# p0 vdd w_587_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_453_311# cin vdd w_506_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1102 a_271_280# p1 vdd w_258_312# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_561_n113# a1 vdd w_548_n81# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 a_381_614# g1 a_424_554# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_883_429# p3p2p1g0 a_883_389# w_877_416# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_693_378# p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 c1 a_445_147# vdd w_504_133# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_304_328# a_271_280# g0 w_291_318# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 a_825_350# p3g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1110 a_564_n389# a3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 s1 a_798_n113# a_876_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_688_664# p1 vdd w_741_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1113 a_797_604# p0 a_797_585# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 vdd a_269_n114# p1 w_258_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1115 p1g0 a_380_291# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_324_n46# b1 a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 a_327_429# a_251_466# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1118 a_693_378# p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 a_380_291# a_304_328# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1120 c2 a_600_239# vdd w_676_271# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 b3 a3 p3 w_368_n380# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1122 a1 b1 a_302_n114# w_328_n116# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 a_328_n37# a_324_n46# a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1124 a_328_97# a_324_88# a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 vdd a3 a_325_n314# w_401_n374# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1126 a_597_n341# a3 b3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 p1p0c0 a_453_311# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1128 a_324_88# b0 a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1129 a_688_664# cin a_797_604# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 vdd g2 a_731_492# w_726_513# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1131 a_883_464# p3p2g1 a_883_429# w_877_451# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_693_378# g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_304_328# p1 g0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1134 g2 a_564_n251# b2 w_584_n213# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1135 a_597_73# a_564_25# b0 w_584_63# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1136 a_597_73# a0 b0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1137 a_771_282# a_738_234# a_816_233# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1138 a_518_635# p1 vdd w_571_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_397_472# g0 vdd w_450_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_797_547# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_496_251# p0 a_496_232# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 a_847_245# a_771_282# vdd w_834_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_597_73# a_564_25# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1147 a_239_604# a_206_556# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1148 a_797_566# p2 a_797_547# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1149 a_453_311# cin a_496_251# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1150 a_453_311# p1 vdd w_440_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 gnd a3 a_325_n314# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1152 a_534_474# p1 vdd w_554_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_304_328# a_271_280# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1154 a_445_147# g0 a_445_140# w_439_134# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 a_797_585# p1 a_797_566# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 gnd a_302_n114# a_269_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_795_n247# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1158 gnd a_269_n114# p1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1159 g0 a_673_36# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1160 a_381_614# g1 vdd w_434_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 s2 c2 a_795_n247# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_561_n113# a1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1163 pocin a_380_153# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_380_153# a_304_190# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1165 a_688_664# p3 vdd w_675_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1166 s3 a_808_n381# a_886_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1167 a_673_n378# a_597_n341# vdd w_660_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 g2 a2 b2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 p1g0 a_380_291# vdd w_400_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1170 c2 a_600_239# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 g1 a_670_n102# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1172 a0 b0 a_302_20# w_328_18# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 a_380_291# a_304_328# vdd w_367_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_688_664# p2 vdd w_708_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1175 p2p1g0 a_397_472# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1176 gnd a2 a_325_n180# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 vdd pocin a_445_140# w_439_167# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1178 c3 a_693_378# vdd w_790_410# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_304_190# p0 cin Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1180 s3 c3 a_808_n381# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1181 a_251_466# a_218_418# g1 w_238_456# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1182 s3 c3 p3 w_867_n335# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 vdd a1 a_324_n46# w_400_n106# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1184 a_673_36# a_597_73# vdd w_660_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1185 a_397_472# g0 a_440_412# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 a_808_n381# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1187 a_798_n113# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_564_25# a0 vdd w_551_57# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 g3 a_673_n378# vdd w_693_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# p2 vdd w_384_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 vdd a_302_n114# a_269_n114# w_291_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1192 a_617_318# p1g0 a_617_278# w_611_305# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1193 a_771_282# cin p0 w_797_280# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 a_738_234# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1195 a_594_n65# a_561_n113# b1 w_581_n75# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_518_635# p2 vdd w_538_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 b0 a0 a_302_20# w_367_22# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_496_232# p1 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1199 a_397_472# p1 vdd w_417_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_206_556# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1201 p3p2p1p0c0 a_688_664# vdd w_845_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 a_610_414# p0 a_610_395# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_534_474# p2 vdd w_521_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_271_142# p0 vdd w_258_174# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1205 s0 a_847_245# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 vdd g1 a_617_318# w_611_340# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 c4 a_825_350# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1208 gnd a1 a_324_n46# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1209 gnd a0 a_324_88# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 gnd a_302_20# a_269_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1211 a_381_614# p2 vdd w_401_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1212 a2 b2 p2 w_329_n250# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 a_251_466# a_218_418# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 a_534_474# cin a_610_414# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1215 a_771_282# cin a_738_234# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 a_381_614# p3 vdd w_368_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1217 p3g2 a_315_567# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1218 a_600_239# g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1219 s2 c2 p2 w_854_n201# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 w_571_625# p1 0.026996f
C1 w_328_n116# a_302_n114# 0.007992f
C2 w_400_n106# a_324_n46# 0.013216f
C3 w_657_n70# a_594_n65# 0.026907f
C4 a_534_474# a_610_414# 0.41238f
C5 a_564_25# vdd 0.439891f
C6 a_302_20# gnd 0.190422f
C7 w_291_318# a_271_280# 0.026794f
C8 a2 a_325_n180# 0.060798f
C9 a_206_556# gnd 0.20619f
C10 p2 c2 0.015947f
C11 w_291_318# vdd 6.13e-19
C12 g2 p2p1p0c0 0.054984f
C13 c1 s1 0.685068f
C14 a_597_73# vdd 0.013824f
C15 w_335_599# vdd 0.008451f
C16 g2 a2 0.012963f
C17 w_867_n335# s3 0.007992f
C18 a_518_635# vdd 1.76176f
C19 p1g0 a_617_278# 0.004158f
C20 a_534_474# p1 0.004034f
C21 w_708_654# a_688_664# 0.027639f
C22 a_600_239# p1p0c0 0.206583f
C23 a_453_311# p0 0.005763f
C24 a_884_498# p3g2 3.63e-19
C25 a_738_234# gnd 0.206673f
C26 cin vdd 0.024447f
C27 w_551_n357# vdd 0.0086f
C28 w_693_n346# a_673_n378# 0.026907f
C29 w_554_464# vdd 0.008451f
C30 a_381_614# p3p2g1 0.060798f
C31 a_594_556# p2 0.013746f
C32 w_877_451# p3p2g1 0.036563f
C33 w_725_444# a_731_417# 0.008113f
C34 w_725_411# p2p1p0c0 0.001174f
C35 p1g0 vdd 0.439883f
C36 a_771_282# gnd 0.190422f
C37 a1 a_302_n114# 0.413834f
C38 w_450_462# g0 0.026794f
C39 w_604_625# a_518_635# 0.027639f
C40 w_401_n374# a3 0.028034f
C41 w_368_n380# b3 0.01395f
C42 w_551_n219# vdd 0.008518f
C43 w_335_599# p3g2 0.013216f
C44 a_424_554# a_424_535# 0.41238f
C45 a_594_556# a_594_537# 0.41238f
C46 w_238_456# vdd 6.13e-19
C47 a_381_614# p2 0.005763f
C48 w_439_167# pocin 0.036563f
C49 w_854_n201# c3 5.29e-20
C50 c4 vdd 0.439883f
C51 w_725_479# p2p1g0 0.036563f
C52 w_878_485# a_883_464# 0.009864f
C53 a_610_377# gnd 0.41238f
C54 a_304_328# a_380_291# 0.060798f
C55 w_657_n70# vdd 0.008507f
C56 w_642_625# vdd 0.008451f
C57 p3 a_424_535# 0.013746f
C58 a_797_585# a_797_566# 0.41238f
C59 g3 vdd 0.442872f
C60 w_620_464# a_534_474# 0.027639f
C61 b0 a_328_97# 0.001802f
C62 a_324_88# a_302_20# 0.286223f
C63 w_488_462# p2p1g0 0.013216f
C64 a_597_73# a_564_25# 0.003752f
C65 w_725_479# a_731_492# 0.01128f
C66 c3 gnd 0.223819f
C67 w_693_68# vdd 0.008451f
C68 w_401_n240# a_325_n180# 0.013216f
C69 a_325_n314# a_329_n305# 0.14502f
C70 w_815_n209# p2 0.028748f
C71 a_518_635# a_594_575# 0.41238f
C72 w_725_266# a_738_234# 0.013216f
C73 a3 a_564_n389# 0.060856f
C74 a_564_n251# gnd 0.20619f
C75 p2p1p0c0 vdd 0.439883f
C76 w_384_462# p2 0.026794f
C77 w_417_462# a_397_472# 0.027639f
C78 a_693_378# gnd 1.08291f
C79 p2 g1 0.127859f
C80 w_258_17# vdd 0.008451f
C81 w_818_n75# s1 0.015055f
C82 w_302_599# a_239_604# 0.026907f
C83 w_867_n335# p3 0.007896f
C84 a_798_n113# gnd 0.206673f
C85 w_611_305# p1g0 0.036782f
C86 w_611_272# a_600_239# 0.013329f
C87 w_544_301# p1p0c0 0.013216f
C88 w_439_167# g0 4.29e-19
C89 a2 vdd 0.195509f
C90 c3 c2 4.66e-20
C91 a_397_472# gnd 0.042086f
C92 w_314_461# a_251_466# 0.026907f
C93 a_218_418# vdd 0.439891f
C94 a_397_472# g0 0.059018f
C95 w_867_277# vdd 0.008451f
C96 p2p1p0c0 a_731_417# 0.004158f
C97 w_581_n75# a_561_n113# 0.026794f
C98 w_657_n70# a_670_n102# 0.013216f
C99 a_693_378# p2g1 0.206583f
C100 a_324_n46# gnd 0.206673f
C101 w_544_301# a_453_311# 0.027163f
C102 w_368_n380# p3 0.015055f
C103 a_797_547# gnd 0.41238f
C104 a_251_466# vdd 0.017997f
C105 p0 a_496_232# 0.013746f
C106 c3 c1 2.14e-19
C107 a_883_464# a_883_429# 0.41238f
C108 w_581_n75# a_594_n65# 0.019526f
C109 w_400_n106# b1 0.015139f
C110 w_548_n81# a1 0.02809f
C111 w_291_n117# a_302_n114# 0.027261f
C112 w_611_340# vdd 0.013119f
C113 w_587_464# p0 0.026996f
C114 a_673_36# vdd 0.441416f
C115 a2 b2 0.531092f
C116 a_269_20# gnd 0.248155f
C117 w_400_323# a_380_291# 0.026907f
C118 w_258_312# a_271_280# 0.013216f
C119 p2 a_329_n171# 0.20619f
C120 a_315_567# gnd 0.248155f
C121 w_258_312# vdd 0.0086f
C122 p1 s1 0.413834f
C123 c1 a_798_n113# 0.016996f
C124 pocin gnd 0.372676f
C125 a_445_140# vdd 0.41238f
C126 w_302_599# vdd 0.008507f
C127 w_675_654# a_688_664# 0.017642f
C128 w_642_625# a_518_635# 0.027163f
C129 p2 p1 2.50865f
C130 a_688_664# vdd 2.20188f
C131 w_828_n343# s3 0.015055f
C132 a_600_239# a_617_278# 0.453641f
C133 w_584_63# b0 0.008938f
C134 w_367_22# a_302_20# 0.015055f
C135 a_304_190# gnd 0.701773f
C136 a_269_n114# p1 0.060798f
C137 p0 vdd 0.678634f
C138 w_584_n351# a_564_n389# 0.026794f
C139 w_660_n346# a_673_n378# 0.013216f
C140 w_401_n374# vdd 0.008451f
C141 a_610_395# p0 0.013746f
C142 a_424_554# p2 0.013746f
C143 w_521_464# vdd 0.008451f
C144 b1 a_324_n46# 0.02927f
C145 a_600_239# vdd 0.001532f
C146 w_725_444# p2p1p0c0 0.036782f
C147 w_329_n384# b3 0.027716f
C148 w_368_n380# a3 0.028748f
C149 w_401_n240# vdd 0.008451f
C150 w_401_604# p2 0.026996f
C151 s3 a_886_n382# 0.20619f
C152 w_400_185# pocin 0.013216f
C153 w_205_450# vdd 0.0086f
C154 p3p2p1p0c0 vdd 0.439883f
C155 w_878_485# p3g2 0.036563f
C156 g0 gnd 0.207724f
C157 w_581_n75# vdd 2.04e-19
C158 w_782_n215# a_795_n247# 0.013216f
C159 w_854_n201# c2 0.027735f
C160 w_226_594# g2 0.018971f
C161 a_564_n389# vdd 0.439891f
C162 w_258_174# p0 0.028034f
C163 a_325_n314# gnd 0.206673f
C164 p3 a_594_537# 0.013746f
C165 a_597_73# a_673_36# 0.060798f
C166 w_878_485# a_884_498# 0.01128f
C167 p2g1 gnd 0.207724f
C168 w_587_464# a_534_474# 0.027639f
C169 b0 a_302_20# 0.685117f
C170 p3p2p1g0 vdd 0.439883f
C171 c3 s3 0.692464f
C172 w_571_625# vdd 0.008451f
C173 w_660_68# vdd 0.008507f
C174 w_401_n240# b2 0.015139f
C175 w_551_n219# a2 0.028079f
C176 w_472_604# a_381_614# 0.027163f
C177 w_505_625# p3 0.026794f
C178 a_597_n341# a_564_n389# 0.003752f
C179 b3 a_329_n305# 0.001802f
C180 w_782_n215# p2 0.028034f
C181 p3 a_206_556# 0.060798f
C182 c2 gnd 0.206382f
C183 w_384_462# a_397_472# 0.017642f
C184 w_238_456# a_218_418# 0.026794f
C185 w_504_133# vdd 0.008451f
C186 w_857_n67# c1 0.027735f
C187 w_193_588# p3 0.028034f
C188 w_226_594# a_239_604# 0.019526f
C189 w_828_n343# p3 0.028748f
C190 c1 gnd 0.206382f
C191 g0 c1 0.008006f
C192 a_534_474# vdd 1.76176f
C193 w_708_654# p2 0.026794f
C194 a_327_429# gnd 0.248155f
C195 w_238_456# a_251_466# 0.019526f
C196 a_610_377# p1 0.013746f
C197 a_688_664# cin 0.059018f
C198 w_548_n81# a_561_n113# 0.013216f
C199 p2 a_440_393# 0.013746f
C200 w_834_277# vdd 0.008507f
C201 w_329_n384# p3 0.007992f
C202 a_302_n114# vdd 0.019283f
C203 b1 gnd 0.035378f
C204 w_506_301# a_453_311# 0.027639f
C205 p0 cin 0.015947f
C206 a_304_190# a_271_142# 0.003752f
C207 w_400_n106# a1 0.028034f
C208 w_291_n117# a_269_n114# 0.013216f
C209 w_367_n112# b1 0.01395f
C210 a_883_464# p3p2g1 3.63e-19
C211 p2p1g0 a_693_378# 0.001345f
C212 a_327_429# p2g1 0.060798f
C213 w_544_301# vdd 0.008451f
C214 w_367_323# a_380_291# 0.013216f
C215 a_324_88# gnd 0.206673f
C216 w_538_625# vdd 0.008451f
C217 p2 a_325_n180# 0.288532f
C218 a_381_614# gnd 0.042086f
C219 w_693_68# a_673_36# 0.026907f
C220 w_942_382# vdd 0.008451f
C221 a_397_472# p2p1g0 0.060798f
C222 p1 a_798_n113# 0.060798f
C223 a_445_147# vdd 0.001532f
C224 a_271_142# gnd 0.20619f
C225 w_226_594# vdd 6.13e-19
C226 a_600_239# p1g0 0.040556f
C227 p3 a_329_n305# 0.20619f
C228 a_397_472# p1 0.005763f
C229 a_518_635# p3p2p1g0 0.060798f
C230 w_328_18# a_302_20# 0.007992f
C231 a_251_466# a_218_418# 0.003752f
C232 p3 c3 0.028649f
C233 w_400_28# a_324_88# 0.013216f
C234 w_660_68# a_597_73# 0.026907f
C235 g2 p2 0.073455f
C236 w_571_625# a_518_635# 0.027639f
C237 s0 vdd 0.439883f
C238 w_790_410# c3 0.013216f
C239 w_551_n357# a_564_n389# 0.013216f
C240 a_797_566# p2 0.013746f
C241 w_488_462# vdd 0.008451f
C242 a_847_245# vdd 0.441416f
C243 a1 a_324_n46# 0.060798f
C244 g1 gnd 0.367778f
C245 w_790_410# a_693_378# 0.027289f
C246 w_329_n384# a3 0.007896f
C247 w_845_654# vdd 0.008451f
C248 a_206_556# g2 0.008991f
C249 w_258_17# p0 0.013216f
C250 a_808_n381# a_886_n382# 0.14502f
C251 a_380_291# vdd 0.441416f
C252 a_304_328# gnd 0.701773f
C253 a_883_389# p3p2p1p0c0 0.015843f
C254 w_548_n81# vdd 0.0086f
C255 a_534_474# cin 0.059018f
C256 w_815_n209# c2 0.01352f
C257 a_304_328# g0 0.753587f
C258 w_193_588# g2 0.009535f
C259 p3 a_797_547# 0.013746f
C260 b3 gnd 0.034146f
C261 w_367_185# a_304_190# 0.026907f
C262 a_673_n378# vdd 0.441416f
C263 c3 a_808_n381# 0.017003f
C264 a_825_350# vdd 0.001532f
C265 w_642_625# p3p2p1g0 0.013216f
C266 w_726_513# a_731_492# 0.009864f
C267 w_554_464# a_534_474# 0.027639f
C268 a0 a_302_20# 0.413834f
C269 p3p2p1g0 a_883_389# 0.004158f
C270 w_401_n240# a2 0.028034f
C271 w_368_n246# b2 0.01395f
C272 w_584_63# vdd 2.04e-19
C273 w_538_625# a_518_635# 0.027639f
C274 w_434_604# a_381_614# 0.027639f
C275 b3 a_325_n314# 0.02927f
C276 a_239_604# a_206_556# 0.003752f
C277 a_795_n247# vdd 0.439891f
C278 w_417_462# p1 0.026996f
C279 a_597_n341# a_673_n378# 0.060798f
C280 w_205_450# a_218_418# 0.013216f
C281 p2p1g0 gnd 0.207724f
C282 p3p2g1 vdd 0.439963f
C283 a_797_585# p0 0.013746f
C284 a_883_429# a_883_389# 0.41238f
C285 w_857_n67# p1 0.007896f
C286 w_818_n75# c1 0.01352f
C287 a_797_604# cin 0.013746f
C288 w_785_n81# a_798_n113# 0.013216f
C289 w_795_n349# p3 0.028034f
C290 s2 a_873_n248# 0.20619f
C291 p1 gnd 0.684683f
C292 w_726_513# p3 4.5e-19
C293 g1 b1 0.281479f
C294 a_380_153# pocin 0.060798f
C295 p2 vdd 0.623899f
C296 w_797_280# vdd 0.001288f
C297 a_688_664# p0 0.005763f
C298 p3g2 a_825_350# 0.001345f
C299 w_473_301# a_453_311# 0.027639f
C300 a1 gnd 1.537765f
C301 a_269_n114# vdd 0.441416f
C302 a_304_190# a_380_153# 0.060798f
C303 w_434_604# g1 0.026794f
C304 a_381_614# g1 0.059018f
C305 a_534_474# p2p1p0c0 0.060798f
C306 w_506_301# vdd 0.008451f
C307 w_258_n117# a_269_n114# 0.026907f
C308 w_328_n116# b1 0.027716f
C309 w_367_n112# a1 0.028748f
C310 a_397_472# a_440_412# 0.41238f
C311 b0 gnd 0.035498f
C312 a_302_20# vdd 0.019283f
C313 w_400_323# g0 0.011382f
C314 w_942_382# c4 0.013216f
C315 w_505_625# vdd 0.008451f
C316 a_206_556# vdd 0.439891f
C317 p2 b2 0.6987f
C318 p3 gnd 1.515037f
C319 g2 a_564_n251# 0.003752f
C320 w_676_271# c2 0.013216f
C321 w_584_63# a_564_25# 0.026794f
C322 w_660_68# a_673_36# 0.013216f
C323 g2 a_693_378# 1.39e-20
C324 a_731_492# a_731_457# 0.41238f
C325 a_688_664# p3p2p1p0c0 0.060798f
C326 a_380_153# gnd 0.248155f
C327 p1 c1 0.015947f
C328 w_193_588# vdd 0.0086f
C329 w_795_n349# a_808_n381# 0.013216f
C330 p3 a_325_n314# 0.286223f
C331 w_584_63# a_597_73# 0.019526f
C332 w_879_518# vdd 0.013167f
C333 w_291_17# a_302_20# 0.027261f
C334 w_400_28# b0 0.015139f
C335 w_551_57# a0 0.028093f
C336 a_738_234# vdd 0.439891f
C337 p1p0c0 gnd 0.207724f
C338 a_302_n114# a_328_n37# 0.20619f
C339 g0 p1p0c0 0.002352f
C340 a_594_556# p1 0.013746f
C341 a_380_291# p1g0 0.060798f
C342 w_450_462# vdd 0.008451f
C343 w_440_301# p1 0.026794f
C344 a1 b1 0.614689f
C345 w_725_411# a_693_378# 0.013329f
C346 a_453_311# gnd 0.042086f
C347 a_771_282# vdd 0.019283f
C348 a_808_n381# gnd 0.206673f
C349 w_400_185# a_380_153# 0.026907f
C350 a_518_635# p2 0.004034f
C351 a_797_566# a_797_547# 0.41238f
C352 w_807_654# vdd 0.008451f
C353 a_440_393# gnd 0.41238f
C354 w_347_461# p2g1 0.013216f
C355 a_534_474# p0 0.005763f
C356 w_400_n106# vdd 0.0086f
C357 w_584_n213# a_564_n251# 0.026794f
C358 a_825_350# c4 0.060798f
C359 a_610_395# a_610_377# 0.41238f
C360 a_673_n378# g3 0.060798f
C361 a_381_614# a_424_554# 0.41238f
C362 w_867_277# s0 0.013216f
C363 a_797_604# a_797_585# 0.41238f
C364 a3 gnd 0.414526f
C365 w_797_280# cin 0.027729f
C366 w_291_180# a_304_190# 0.019526f
C367 w_726_513# g2 0.036563f
C368 a_825_350# g3 1.39e-20
C369 w_521_464# a_534_474# 0.017642f
C370 c3 vdd 0.446487f
C371 b0 a_324_88# 0.02927f
C372 w_879_518# a_884_498# 0.009864f
C373 a_440_412# g0 0.013746f
C374 a_825_350# a_883_389# 0.453641f
C375 w_329_n250# b2 0.027716f
C376 w_368_n246# a2 0.028748f
C377 w_551_57# vdd 0.0086f
C378 w_401_604# a_381_614# 0.027639f
C379 w_505_625# a_518_635# 0.017642f
C380 w_506_301# cin 0.026794f
C381 a_325_n180# gnd 0.206673f
C382 a3 a_325_n314# 0.060798f
C383 a_564_n251# vdd 0.439891f
C384 a_239_604# a_315_567# 0.060798f
C385 p3 a_381_614# 0.002444f
C386 w_867_277# a_847_245# 0.026907f
C387 a_688_664# a_797_604# 0.41238f
C388 a_693_378# vdd 0.001532f
C389 a_445_147# a_445_140# 0.453641f
C390 w_347_461# a_327_429# 0.026907f
C391 w_439_167# vdd 0.010186f
C392 a_883_429# p3p2p1g0 4.37e-21
C393 w_818_n75# p1 0.028748f
C394 a_797_604# p0 0.013746f
C395 a_798_n113# vdd 0.439891f
C396 a_795_n247# a_873_n248# 0.14502f
C397 a_561_n113# gnd 0.20619f
C398 w_741_654# p1 0.026794f
C399 g1 a1 0.115698f
C400 a_304_328# p1 0.001371f
C401 a_397_472# vdd 1.32165f
C402 g2 gnd 0.829522f
C403 cin a_816_233# 0.002154f
C404 w_758_272# vdd 6.13e-19
C405 a_424_554# g1 0.013746f
C406 a_693_378# a_731_417# 0.453641f
C407 a_324_n46# vdd 0.439891f
C408 b2 a_564_n251# 0.002958f
C409 w_440_301# a_453_311# 0.017642f
C410 a_594_n65# gnd 0.701773f
C411 a_738_234# cin 0.017003f
C412 w_328_n116# a1 0.007896f
C413 w_473_301# vdd 0.008451f
C414 p3 g1 0.652627f
C415 w_367_323# g0 0.011382f
C416 a0 gnd 1.211792f
C417 a_269_20# vdd 0.441416f
C418 w_472_604# vdd 0.008451f
C419 w_845_654# a_688_664# 0.027163f
C420 a_771_282# cin 0.685096f
C421 p3 s3 0.413834f
C422 a_315_567# vdd 0.441416f
C423 a_239_604# gnd 0.248155f
C424 p2 a2 0.49284f
C425 a_731_492# p2p1g0 3.63e-19
C426 p2 a_218_418# 0.060798f
C427 w_551_57# a_564_25# 0.013216f
C428 a_496_232# gnd 0.41238f
C429 w_877_383# a_883_389# 0.017071f
C430 pocin vdd 0.439883f
C431 w_807_654# cin 0.026794f
C432 w_795_n349# vdd 0.008518f
C433 a_453_311# a_496_251# 0.41238f
C434 p3 b3 0.685112f
C435 a_617_318# a_617_278# 0.41238f
C436 w_291_17# a_269_20# 0.013216f
C437 w_400_28# a0 0.028034f
C438 w_367_22# b0 0.01395f
C439 w_879_518# g3 0.036563f
C440 w_726_513# vdd 0.013119f
C441 a_251_466# p2 0.001371f
C442 b1 a_561_n113# 0.00343f
C443 w_725_411# p2g1 0.043313f
C444 a_304_190# vdd 0.017997f
C445 c3 cin 5.1e-19
C446 a_315_567# p3g2 0.060798f
C447 w_417_462# vdd 0.008451f
C448 w_504_133# a_445_147# 0.027289f
C449 w_439_134# a_445_140# 0.017071f
C450 a_617_318# vdd 0.41238f
C451 a_271_280# gnd 0.20619f
C452 w_845_654# p3p2p1p0c0 0.013216f
C453 a_594_n65# b1 0.7623f
C454 w_877_451# a_883_464# 0.01128f
C455 g0 a_271_280# 0.001372f
C456 a_808_n381# s3 0.286223f
C457 w_774_654# vdd 0.008451f
C458 a_688_664# p2 0.004034f
C459 w_291_180# a_271_142# 0.026794f
C460 w_367_185# a_380_153# 0.013216f
C461 vdd gnd 2.215758f
C462 g0 vdd 0.56271f
C463 w_367_n112# vdd 6.13e-19
C464 w_551_n219# a_564_n251# 0.013216f
C465 a_825_350# p3p2p1p0c0 0.206583f
C466 w_797_280# p0 0.007896f
C467 w_758_272# cin 0.01352f
C468 a_325_n314# vdd 0.439883f
C469 a_597_n341# gnd 0.701773f
C470 w_521_464# p2 0.026794f
C471 a0 a_324_88# 0.060798f
C472 c3 g3 0.055169f
C473 p2g1 vdd 0.439883f
C474 a_825_350# p3p2p1g0 0.040556f
C475 w_329_n250# a2 0.007896f
C476 w_400_28# vdd 0.0086f
C477 w_368_604# a_381_614# 0.017642f
C478 w_335_599# a_315_567# 0.026907f
C479 w_401_n240# p2 0.003504f
C480 a3 b3 0.535308f
C481 w_834_277# a_847_245# 0.013216f
C482 c2 vdd 0.439883f
C483 b2 gnd 0.037864f
C484 w_604_625# g0 0.026794f
C485 a_453_311# p1 0.002444f
C486 w_205_450# p2 0.028034f
C487 p3g2 gnd 0.207724f
C488 w_314_461# a_327_429# 0.013216f
C489 c3 a_873_n248# 4.29e-20
C490 a_731_417# p2g1 0.015843f
C491 p3p2g1 p3p2p1g0 0.041485f
C492 w_785_n81# p1 0.028034f
C493 w_400_185# vdd 0.008451f
C494 g2 g1 1.63579f
C495 a_795_n247# s2 0.286223f
C496 w_611_305# a_617_318# 0.009864f
C497 c1 vdd 0.439883f
C498 a_670_n102# gnd 0.248155f
C499 a_327_429# vdd 0.441416f
C500 a_440_393# p1 0.013746f
C501 w_725_266# vdd 0.0086f
C502 a_693_378# p2p1p0c0 0.040556f
C503 a_731_457# a_731_417# 0.41238f
C504 w_867_277# c3 3.18e-20
C505 a_564_25# gnd 0.20619f
C506 b1 vdd 0.015576f
C507 a2 a_564_n251# 0.060856f
C508 a_325_n180# a_329_n171# 0.14502f
C509 a_738_234# p0 0.060798f
C510 a_304_190# cin 0.740337f
C511 a_496_251# a_496_232# 0.41238f
C512 p2 s2 0.413834f
C513 a_440_412# p1 0.013746f
C514 g2 b3 3.99e-19
C515 w_440_301# vdd 0.008451f
C516 a_594_575# g0 0.013746f
C517 a_597_73# gnd 0.248155f
C518 w_367_323# a_304_328# 0.026907f
C519 s1 a_876_n114# 0.20619f
C520 a_324_88# vdd 0.439891f
C521 w_877_383# p3p2p1p0c0 0.043313f
C522 w_291_318# g0 0.008451f
C523 w_434_604# vdd 0.008451f
C524 a_381_614# vdd 1.32165f
C525 a_847_245# s0 0.060798f
C526 a_518_635# gnd 0.042086f
C527 w_807_654# a_688_664# 0.027639f
C528 a_771_282# p0 0.413834f
C529 p3 a_808_n381# 0.060798f
C530 a_518_635# g0 0.059018f
C531 p2 a_534_474# 0.002444f
C532 w_942_382# a_825_350# 0.027289f
C533 w_877_416# a_883_389# 0.008113f
C534 w_877_383# p3p2p1g0 0.001142f
C535 cin gnd 1.92e-19
C536 a_271_142# vdd 0.439891f
C537 a_617_318# p1g0 4.37e-21
C538 a_453_311# p1p0c0 0.060798f
C539 w_693_n346# vdd 0.008451f
C540 p3 a3 0.413834f
C541 a_424_535# p2 0.013746f
C542 w_258_17# a_269_20# 0.026907f
C543 w_658_464# vdd 0.008451f
C544 w_328_18# b0 0.027757f
C545 w_367_22# a0 0.028748f
C546 a_269_n114# a_302_n114# 0.060798f
C547 p1g0 gnd 0.207724f
C548 a_324_n46# a_328_n37# 0.14502f
C549 a1 a_561_n113# 0.060856f
C550 c3 p0 1.64e-20
C551 a_797_566# p1 0.013746f
C552 w_584_n351# b3 0.008451f
C553 g0 p1g0 0.007385f
C554 w_538_625# p2 0.026794f
C555 w_690_n70# g1 0.01323f
C556 w_439_167# a_445_140# 0.008113f
C557 w_439_134# a_445_147# 0.013329f
C558 w_384_462# vdd 0.008451f
C559 w_725_444# a_731_457# 0.009864f
C560 c4 gnd 0.20619f
C561 a_594_n65# a1 0.001371f
C562 g1 vdd 0.727672f
C563 a_304_328# a_271_280# 0.003752f
C564 w_258_174# a_271_142# 0.013216f
C565 a_594_575# a_594_556# 0.41238f
C566 g3 gnd 0.207724f
C567 w_741_654# vdd 0.008451f
C568 p3 g2 0.016679f
C569 a_304_328# vdd 0.017767f
C570 a_302_20# a_328_97# 0.20619f
C571 a_496_232# p1 0.013746f
C572 w_328_n116# vdd 0.001288f
C573 w_758_272# p0 0.028748f
C574 w_693_68# g0 0.01325f
C575 b3 vdd 0.013251f
C576 p2p1p0c0 gnd 0.207724f
C577 a0 b0 0.539271f
C578 g1 b2 7.83e-19
C579 w_367_22# vdd 6.13e-19
C580 a_610_414# a_610_395# 0.41238f
C581 a_440_412# a_440_393# 0.41238f
C582 w_368_604# p3 0.026794f
C583 w_302_599# a_315_567# 0.013216f
C584 w_226_594# a_206_556# 0.026794f
C585 w_611_272# p1p0c0 0.043313f
C586 w_473_301# p0 0.026996f
C587 w_368_n246# p2 0.018553f
C588 a_597_n341# b3 0.756931f
C589 a_239_604# p3 0.001371f
C590 a2 gnd 1.559369f
C591 w_834_277# a_771_282# 0.027261f
C592 a_218_418# gnd 0.20619f
C593 pocin a_445_140# 0.185571f
C594 a_271_280# p1 0.060798f
C595 c3 s2 0.015855f
C596 p2p1g0 vdd 0.439883f
C597 p0 a_269_20# 0.060798f
C598 g1 a_670_n102# 0.060798f
C599 p3p2g1 a_825_350# 0.001345f
C600 w_367_185# vdd 0.008507f
C601 w_611_340# a_617_318# 0.009864f
C602 c2 a_873_n248# 0.001866f
C603 p1 vdd 0.649086f
C604 cin a_271_142# 0.001372f
C605 a_731_492# vdd 0.41238f
C606 c3 a_876_n114# 6.44e-19
C607 a_610_395# p1 0.013746f
C608 a_251_466# gnd 0.701773f
C609 w_676_271# vdd 0.008451f
C610 w_611_340# gnd 1.17e-19
C611 a_731_457# p2p1p0c0 4.37e-21
C612 w_258_n117# p1 0.013216f
C613 w_834_277# c3 3.18e-20
C614 a_673_36# gnd 0.248155f
C615 b2 a_329_n171# 0.001802f
C616 a1 vdd 0.229007f
C617 g2 a3 0.009821f
C618 g0 a_673_36# 0.060812f
C619 a_304_190# p0 0.001371f
C620 a_496_251# cin 0.013746f
C621 p2 a_795_n247# 0.060798f
C622 w_400_323# vdd 0.008451f
C623 w_291_318# a_304_328# 0.019526f
C624 b0 vdd 0.015588f
C625 a_798_n113# a_876_n114# 0.14502f
C626 w_401_604# vdd 0.008451f
C627 w_675_654# p3 0.026794f
C628 a_688_664# gnd 0.042086f
C629 a_617_278# p1p0c0 0.015843f
C630 g0 a_445_140# 0.016231f
C631 w_774_654# a_688_664# 0.027639f
C632 p3 vdd 0.976896f
C633 w_790_410# vdd 0.008451f
C634 a_380_153# vdd 0.441416f
C635 w_877_416# p3p2p1g0 0.036782f
C636 w_877_383# a_825_350# 0.013329f
C637 w_774_654# p0 0.026996f
C638 p0 gnd 0.628007f
C639 w_693_n346# g3 0.013222f
C640 a_771_282# a_847_245# 0.060798f
C641 g1 p1g0 0.035992f
C642 w_660_n346# vdd 0.008507f
C643 w_620_464# vdd 0.008451f
C644 w_867_n335# c3 0.027759f
C645 w_328_18# a0 0.007896f
C646 a_594_537# p2 0.013746f
C647 a_251_466# a_327_429# 0.060798f
C648 b1 a_328_n37# 0.001802f
C649 a_594_n65# a_561_n113# 0.003752f
C650 w_877_416# a_883_429# 0.009864f
C651 w_238_456# g1 0.021496f
C652 p1p0c0 vdd 0.439883f
C653 a_324_n46# a_302_n114# 0.286223f
C654 a_600_239# gnd 0.829424f
C655 w_660_n346# a_597_n341# 0.026907f
C656 w_401_n374# a_325_n314# 0.013216f
C657 a_610_414# cin 0.013746f
C658 a_594_575# p1 0.013746f
C659 w_782_n215# vdd 0.008518f
C660 c3 s0 0.003003f
C661 w_347_461# vdd 0.008451f
C662 w_658_464# p2p1p0c0 0.013216f
C663 a_453_311# vdd 1.32165f
C664 p3p2p1p0c0 gnd 0.207724f
C665 c3 a_847_245# 0.006337f
C666 w_785_n81# vdd 0.008518f
C667 w_854_n201# s2 0.007992f
C668 a_518_635# p1 0.005763f
C669 a_239_604# g2 0.75303f
C670 w_708_654# vdd 0.008451f
C671 a_564_n389# gnd 0.20619f
C672 vdd a_808_n381# 0.439891f
C673 a_600_239# c2 0.060798f
C674 p3p2p1g0 gnd 0.207724f
C675 b0 a_564_25# 0.00288f
C676 w_291_n117# vdd 0.008507f
C677 w_725_266# p0 0.028034f
C678 w_554_464# p1 0.026794f
C679 a3 vdd 0.20154f
C680 w_488_462# a_397_472# 0.027163f
C681 a_597_73# b0 0.756776f
C682 g1 a2 0.011016f
C683 c3 a_825_350# 2.29e-19
C684 w_328_18# vdd 0.001288f
C685 a_218_418# g1 0.012164f
C686 w_193_588# a_206_556# 0.013216f
C687 a_597_n341# a3 0.001371f
C688 a_325_n180# vdd 0.439883f
C689 w_797_280# a_771_282# 0.007992f
C690 w_611_272# a_617_278# 0.017071f
C691 w_584_n213# g2 0.019526f
C692 w_504_133# g0 0.011197f
C693 a_518_635# p3 0.002444f
C694 w_329_n250# p2 0.011491f
C695 a_534_474# gnd 0.042086f
C696 pocin a_445_147# 1.39e-20
C697 c3 a_795_n247# 4.01e-19
C698 a_251_466# g1 0.756678f
C699 w_291_180# vdd 6.13e-19
C700 p2 a_610_377# 0.013746f
C701 a_561_n113# vdd 0.439891f
C702 a_302_n114# gnd 0.190422f
C703 w_611_340# g1 0.036563f
C704 w_400_323# p1g0 0.013216f
C705 c2 s2 0.685083f
C706 a_424_535# gnd 0.41238f
C707 p0 a_271_142# 0.060798f
C708 g2 vdd 0.029171f
C709 a_738_234# a_816_233# 0.14502f
C710 c3 s1 0.003481f
C711 p2p1g0 p2p1p0c0 0.041485f
C712 w_581_n75# b1 0.009938f
C713 w_367_n112# a_302_n114# 0.015055f
C714 w_797_280# c3 0.013839f
C715 b2 a_325_n180# 0.02927f
C716 a_594_n65# vdd 0.013824f
C717 w_620_464# cin 0.026794f
C718 w_544_301# g0 0.00229f
C719 a_496_251# p0 0.013746f
C720 a_771_282# a_816_233# 0.20619f
C721 p2 a_564_n251# 0.002692f
C722 g2 a_597_n341# 0.013288f
C723 w_504_133# c1 0.013216f
C724 w_367_323# vdd 0.008493f
C725 a_798_n113# s1 0.286223f
C726 a_445_147# gnd 0.575941f
C727 a0 vdd 0.234154f
C728 c1 a_876_n114# 0.001856f
C729 w_368_604# vdd 0.008451f
C730 a_771_282# a_738_234# 0.286223f
C731 g0 a_445_147# 0.216537f
C732 w_741_654# a_688_664# 0.027639f
C733 a_453_311# cin 0.059018f
C734 g2 b2 0.764942f
C735 a_239_604# vdd 0.017997f
C736 a_397_472# p2 0.002444f
C737 a_884_498# a_883_464# 0.41238f
C738 s0 gnd 0.20619f
C739 g1 a_600_239# 1.39e-20
C740 w_472_604# p3p2g1 0.013216f
C741 w_587_464# vdd 0.008451f
C742 a_797_547# p2 0.013746f
C743 w_828_n343# c3 0.016729f
C744 a_847_245# gnd 0.248155f
C745 b1 a_302_n114# 0.685112f
C746 w_205_450# g1 0.013044f
C747 w_725_411# a_731_417# 0.017071f
C748 w_877_451# a_883_429# 0.009864f
C749 a_594_n65# a_670_n102# 0.060798f
C750 a_797_585# p1 0.013746f
C751 w_401_n374# b3 0.015139f
C752 w_551_n357# a3 0.02808f
C753 w_584_n351# a_597_n341# 0.019526f
C754 a_610_414# p0 0.013746f
C755 w_439_134# pocin 1.21e-19
C756 w_258_312# p1 0.028034f
C757 w_314_461# vdd 0.008507f
C758 a_271_280# vdd 0.439891f
C759 w_725_479# a_731_457# 0.009864f
C760 a_445_147# c1 0.060798f
C761 a_380_291# gnd 0.248155f
C762 w_690_n70# vdd 0.008451f
C763 w_815_n209# s2 0.015055f
C764 g0 a_380_291# 0.008577f
C765 c3 a_771_282# 0.008546f
C766 a_688_664# p1 0.004034f
C767 w_675_654# vdd 0.008451f
C768 a_673_n378# gnd 0.248155f
C769 w_291_180# cin 0.008451f
C770 a0 a_564_25# 0.060867f
C771 c3 a_886_n382# 0.002154f
C772 a_269_20# a_302_20# 0.060798f
C773 a_825_350# gnd 1.35993f
C774 w_658_464# a_534_474# 0.027163f
C775 a_324_88# a_328_97# 0.14502f
C776 w_584_n213# b2 0.008451f
C777 w_258_n117# vdd 0.008451f
C778 a_597_n341# vdd 0.011738f
C779 b3 a_564_n389# 0.00288f
C780 a_795_n247# gnd 0.206673f
C781 w_854_n201# p2 0.007896f
C782 w_450_462# a_397_472# 0.027639f
C783 p3p2g1 gnd 0.207724f
C784 a_597_73# a0 0.001371f
C785 w_291_17# vdd 0.008507f
C786 w_857_n67# s1 0.007992f
C787 w_604_625# vdd 0.008451f
C788 w_439_134# g0 0.051057f
C789 w_758_272# a_771_282# 0.015055f
C790 a_688_664# p3 0.002444f
C791 w_611_305# a_617_278# 0.008113f
C792 w_611_272# p1g0 0.001158f
C793 w_676_271# a_600_239# 0.027289f
C794 b2 vdd 2.33e-19
C795 p3g2 vdd 0.440124f
C796 p2 gnd 1.655567f
C797 w_690_n70# a_670_n102# 0.026907f
C798 a_693_378# c3 0.060798f
C799 w_258_174# vdd 0.0086f
C800 p2 g0 0.0099f
C801 c2 a_795_n247# 0.017003f
C802 a_670_n102# vdd 0.441416f
C803 a_269_n114# gnd 0.248155f
C804 c3 a_798_n113# 0.001329f
C805 a_594_537# gnd 0.41238f
C806 a_884_498# vdd 0.41238f
C807 a_886_n382# 0 0.016528f  
C808 gnd 0 15.638858f  
C809 s3 0 0.473154f  
C810 a_808_n381# 0 0.526842f  
C811 vdd 0 26.588215f  
C812 g3 0 1.71886f  
C813 a_564_n389# 0 0.477455f  
C814 a_673_n378# 0 0.382299f  
C815 a_329_n305# 0 0.016528f  
C816 a_325_n314# 0 0.526842f  
C817 b3 0 6.62907f  
C818 a3 0 2.45012f  
C819 a_597_n341# 0 0.771781f  
C820 a_873_n248# 0 0.016528f  
C821 s2 0 0.462937f  
C822 a_795_n247# 0 0.526842f  
C823 a_564_n251# 0 0.477455f  
C824 c2 0 1.69805f  
C825 a_329_n171# 0 0.016528f  
C826 a_325_n180# 0 0.526842f  
C827 b2 0 6.55321f  
C828 a2 0 2.34823f  
C829 a_876_n114# 0 0.016528f  
C830 s1 0 0.462937f  
C831 a_798_n113# 0 0.526842f  
C832 c1 0 1.7056f  
C833 p1 0 6.214168f  
C834 a_561_n113# 0 0.477455f  
C835 a_670_n102# 0 0.382299f  
C836 a_328_n37# 0 0.016528f  
C837 a_302_n114# 0 0.662497f  
C838 a_269_n114# 0 0.382299f  
C839 a_324_n46# 0 0.526842f  
C840 b1 0 5.6743f  
C841 a1 0 2.37347f  
C842 a_594_n65# 0 0.771781f  
C843 a_564_25# 0 0.477455f  
C844 a_673_36# 0 0.382299f  
C845 a_328_97# 0 0.016528f  
C846 a_302_20# 0 0.662497f  
C847 a_269_20# 0 0.382299f  
C848 a_324_88# 0 0.526842f  
C849 b0 0 6.55448f  
C850 a0 0 2.49553f  
C851 a_597_73# 0 0.804448f  
C852 a_445_140# 0 0.179875f  
C853 a_445_147# 0 1.02677f  
C854 a_816_233# 0 0.016528f  
C855 pocin 0 0.600283f  
C856 a_271_142# 0 0.477455f  
C857 a_380_153# 0 0.382299f  
C858 a_496_232# 0 0.040245f  
C859 cin 0 3.07338f  
C860 p0 0 3.844454f  
C861 s0 0 0.145867f  
C862 a_738_234# 0 0.526842f  
C863 a_304_190# 0 0.771781f  
C864 a_496_251# 0 0.040245f  
C865 p1p0c0 0 0.361176f  
C866 a_617_278# 0 0.206277f  
C867 p1g0 0 1.282447f  
C868 a_600_239# 0 1.28245f  
C869 a_847_245# 0 0.382299f  
C870 a_771_282# 0 0.662497f  
C871 a_617_318# 0 0.150155f  
C872 g1 0 12.668234f  
C873 a_453_311# 0 1.70512f  
C874 a_271_280# 0 0.477455f  
C875 c4 0 0.15567f  
C876 p3p2p1p0c0 0 0.361176f  
C877 a_380_291# 0 0.382299f  
C878 a_610_377# 0 0.036687f  
C879 g0 0 11.042208f  
C880 a_304_328# 0 0.771781f  
C881 a_440_393# 0 0.040245f  
C882 a_610_395# 0 0.040245f  
C883 a_883_389# 0 0.206277f  
C884 p3p2p1g0 0 1.29225f  
C885 a_825_350# 0 1.81546f  
C886 c3 0 2.78154f  
C887 p2g1 0 0.351373f  
C888 a_610_414# 0 0.040245f  
C889 a_440_412# 0 0.040245f  
C890 a_731_417# 0 0.206277f  
C891 p2p1p0c0 0 1.29452f  
C892 a_883_429# 0 0.150155f  
C893 p3p2g1 0 0.681984f  
C894 a_693_378# 0 1.55643f  
C895 a_731_457# 0 0.150155f  
C896 p2p1g0 0 0.681984f  
C897 a_883_464# 0 0.148414f  
C898 p3g2 0 0.859094f  
C899 a_218_418# 0 0.477455f  
C900 a_534_474# 0 2.1423f  
C901 p2 0 8.949098f  
C902 a_397_472# 0 1.70512f  
C903 a_327_429# 0 0.382299f  
C904 a_731_492# 0 0.148414f  
C905 g2 0 17.347467f  
C906 a_884_498# 0 0.144831f  
C907 a_251_466# 0 0.770807f  
C908 a_424_535# 0 0.040245f  
C909 a_594_537# 0 0.040245f  
C910 a_797_547# 0 0.040245f  
C911 a_594_556# 0 0.040245f  
C912 a_424_554# 0 0.040245f  
C913 a_797_566# 0 0.040245f  
C914 a_594_575# 0 0.040245f  
C915 a_797_585# 0 0.040245f  
C916 a_797_604# 0 0.040245f  
C917 a_206_556# 0 0.477455f  
C918 a_315_567# 0 0.382299f  
C919 a_381_614# 0 1.70512f  
C920 p3 0 9.529533f  
C921 a_239_604# 0 0.804448f  
C922 a_518_635# 0 2.1423f  
C923 a_688_664# 0 2.57948f  
C924 w_867_n335# 0 1.25349f  
C925 w_828_n343# 0 1.34991f  
C926 w_795_n349# 0 1.34991f  
C927 w_693_n346# 0 1.34991f  
C928 w_660_n346# 0 1.34991f  
C929 w_584_n351# 0 1.34991f  
C930 w_551_n357# 0 1.34991f  
C931 w_401_n374# 0 1.34991f  
C932 w_368_n380# 0 1.34991f  
C933 w_329_n384# 0 1.25349f  
C934 w_854_n201# 0 1.25349f  
C935 w_815_n209# 0 1.34991f  
C936 w_782_n215# 0 1.34991f  
C937 w_584_n213# 0 1.34991f  
C938 w_551_n219# 0 1.34991f  
C939 w_401_n240# 0 1.34991f  
C940 w_368_n246# 0 1.34991f  
C941 w_329_n250# 0 1.25349f  
C942 w_857_n67# 0 1.25349f  
C943 w_818_n75# 0 1.34991f  
C944 w_785_n81# 0 1.34991f  
C945 w_690_n70# 0 1.34991f  
C946 w_657_n70# 0 1.34991f  
C947 w_581_n75# 0 1.34991f  
C948 w_548_n81# 0 1.34991f  
C949 w_400_n106# 0 1.34991f  
C950 w_367_n112# 0 1.34991f  
C951 w_328_n116# 0 1.25349f  
C952 w_291_n117# 0 1.34991f  
C953 w_258_n117# 0 1.34991f  
C954 w_693_68# 0 1.34991f  
C955 w_660_68# 0 1.34991f  
C956 w_584_63# 0 1.34991f  
C957 w_551_57# 0 1.34991f  
C958 w_400_28# 0 1.34991f  
C959 w_367_22# 0 1.34991f  
C960 w_328_18# 0 1.25349f  
C961 w_291_17# 0 1.34991f  
C962 w_258_17# 0 1.34991f  
C963 w_504_133# 0 1.34991f  
C964 w_439_134# 0 1.34991f  
C965 w_439_167# 0 1.34991f  
C966 w_400_185# 0 1.34991f  
C967 w_367_185# 0 1.34991f  
C968 w_291_180# 0 1.34991f  
C969 w_258_174# 0 1.34991f  
C970 w_867_277# 0 1.34991f  
C971 w_834_277# 0 1.34991f  
C972 w_797_280# 0 1.25349f  
C973 w_758_272# 0 1.34991f  
C974 w_725_266# 0 1.34991f  
C975 w_676_271# 0 1.34991f  
C976 w_611_272# 0 1.34991f  
C977 w_611_305# 0 1.34991f  
C978 w_611_340# 0 1.34991f  
C979 w_544_301# 0 1.34991f  
C980 w_506_301# 0 1.34991f  
C981 w_473_301# 0 1.34991f  
C982 w_440_301# 0 1.34991f  
C983 w_400_323# 0 1.34991f  
C984 w_367_323# 0 1.34991f  
C985 w_291_318# 0 1.34991f  
C986 w_258_312# 0 1.34991f  
C987 w_942_382# 0 1.34991f  
C988 w_877_383# 0 1.34991f  
C989 w_877_416# 0 1.34991f  
C990 w_877_451# 0 1.34991f  
C991 w_790_410# 0 1.34991f  
C992 w_725_411# 0 1.34991f  
C993 w_725_444# 0 1.34991f  
C994 w_878_485# 0 1.34991f  
C995 w_725_479# 0 1.34991f  
C996 w_879_518# 0 1.34991f  
C997 w_726_513# 0 1.34991f  
C998 w_658_464# 0 1.34991f  
C999 w_620_464# 0 1.34991f  
C1000 w_587_464# 0 1.34991f  
C1001 w_554_464# 0 1.34991f  
C1002 w_521_464# 0 1.34991f  
C1003 w_488_462# 0 1.34991f  
C1004 w_450_462# 0 1.34991f  
C1005 w_417_462# 0 1.34991f  
C1006 w_384_462# 0 1.34991f  
C1007 w_347_461# 0 1.34991f  
C1008 w_314_461# 0 1.34991f  
C1009 w_238_456# 0 1.34991f  
C1010 w_205_450# 0 1.34991f  
C1011 w_845_654# 0 1.34991f  
C1012 w_807_654# 0 1.34991f  
C1013 w_774_654# 0 1.34991f  
C1014 w_741_654# 0 1.34991f  
C1015 w_708_654# 0 1.34991f  
C1016 w_675_654# 0 1.34991f  
C1017 w_642_625# 0 1.34991f  
C1018 w_604_625# 0 1.34991f  
C1019 w_571_625# 0 1.34991f  
C1020 w_538_625# 0 1.34991f  
C1021 w_505_625# 0 1.34991f  
C1022 w_472_604# 0 1.34991f  
C1023 w_434_604# 0 1.34991f  
C1024 w_401_604# 0 1.34991f  
C1025 w_368_604# 0 1.34991f  
C1026 w_335_599# 0 1.34991f  
C1027 w_302_599# 0 1.34991f  
C1028 w_226_594# 0 1.34991f  
C1029 w_193_588# 0 1.34991f  




 

* * RISING AND FALLING DELAY MEASUREMENT
* * * Measure the delay for the final carry-out signal (C4)
.measure tran delay_C4_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(c4) VAL=0.9 FALL=1
.measure tran delay_C4_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(c4) VAL=0.9 RISE=1

* * Measure the delay for each sum signal
.measure tran delay_S0_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s0) VAL=0.9 FALL=1
.measure tran delay_S0_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s0) VAL=0.9 RISE=1
.measure tran delay_S1_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s1) VAL=0.9 FALL=1
.measure tran delay_S1_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s1) VAL=0.9 RISE=1
.measure tran delay_S2_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s2) VAL=0.9 FALL=1
.measure tran delay_S2_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s2) VAL=0.9 RISE=1
.measure tran delay_S3_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s3) VAL=0.9 FALL=1
.measure tran delay_S3_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s3) VAL=0.9 RISE=1



.control
  set hcopypscolor = 1             
  set color0 = white               
  set color1 = black               
  set color2 = red                 
  set color3 = blue                
  set color4 = coral               
  set color5 = brown    
  set color6 = cyan
  set color7 = chocolate   
  set color8 = chocolate
  set color9 = blueviolet
  set color10 = cadetblue        
  * for testing        
  * tran 1n 160n
  * for delay  
  tran 0.01n 40n 
   plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+g0 20+g1 22+g2 24+g3   
  plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+p0 20+p1 22+p2 24+p3                      
  * plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+s0 20+s1 22+s2 24+s3                      
    plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+c4 20+s0 22+s1 24+s2 26+s3   
    plot pocin 2+g0 4+c1
    * plot g3 2+p3g2 4+p3p2g1 6+p3p2p1g0 8+p3p2p1p0c0 10+c4 
    plot c1 2+p1 4+s1
  plot s0 2+s1 4+s2 6+s3    
        
.endc