* SPICE3 file created from and.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* Test Signals
Vclk b gnd PULSE(0 'SUPPLY' 0 0.001n 0.01n 10n 20n)
Vd a gnd PULSE(0 'SUPPLY' 0n 0.001n 0.01n 35n 70n)



M1000 y-d abar gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 ybar y-d gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 y ybar vdd w_126_9# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1003 y-d a b Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1004 abar a gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 ybar y-d vdd w_93_9# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 y-d abar b w_17_4# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 abar a vdd w_n16_n2# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 y ybar gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
C0 y-d w_17_4# 2.82f
C1 y-d vdd 1.89f
C2 w_17_4# abar 1.014f
C3 y-d w_93_9# 1.014f
C4 w_n16_n2# vdd 1.128f
C5 ybar w_126_9# 1.014f
C6 a w_n16_n2# 1.014f
C7 vdd w_126_9# 1.128f
C8 y w_126_9# 1.88f
C9 w_93_9# ybar 1.88f
C10 w_17_4# b 1.128f
C11 w_93_9# vdd 1.128f
C12 w_n16_n2# abar 1.88f
C13 b vdd 1.26f
C14 gnd 0 77.456f 
C15 y 0 3.76f 
C16 vdd 0 38.429f 
C17 abar 0 18.082f 
C18 ybar 0 14.266f 
C19 b 0 8.177999f 
C20 a 0 44.896f 
C21 y-d 0 44.863f 


.control
  set hcopypscolor = 1
  set color0 = white
  set color1 = black
  set color2 = red
  set color3 = blue
  set color4 = brown
  set color5 = magenta
  set color6 = cyan
  set color7 = green
  tran 1n 200n
    plot a 2+b 4+y
.endc
