* Positive-Edge-Triggered D Flip-Flop - TSPS Design 
* TSMC 180nm Technology Parameters
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* Test Signals
Vclk clk gnd PULSE(0 'SUPPLY' 0 1n 1n 10n 20n)
Vd d gnd PULSE(0 'SUPPLY' 10n 1n 1n 10n 40n)




* SPICE3 file created from dff.ext - technology: scmos

.option scale=90n

M1000 a_n214_n85# d gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 vdd d a_n206_n60# w_n216_n43# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1002 q qbar vdd w_n23_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1003 a_n82_n85# a_n137_n36# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1004 qbar clk a_n82_n85# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 a_n144_n85# clk gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1006 a_n206_n60# clk a_n214_n85# w_n216_n73# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 vdd a_n137_n36# qbar w_n85_n43# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 a_n137_n36# a_n214_n85# a_n144_n85# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1009 q qbar gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1010 vdd clk a_n137_n36# w_n147_n43# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 clk a_n144_n85# 0.011946f
C1 a_n137_n36# a_n214_n85# 4.83e-19
C2 w_n216_n73# a_n206_n60# 0.006024f
C3 qbar vdd 0.413752f
C4 w_n147_n43# a_n137_n36# 0.0075f
C5 clk a_n82_n85# 1.92e-20
C6 a_n137_n36# a_n144_n85# 0.20619f
C7 d gnd 7.27e-19
C8 w_n85_n43# a_n137_n36# 0.028451f
C9 w_n216_n73# clk 0.041363f
C10 a_n137_n36# a_n82_n85# 0.096222f
C11 vdd d 7.27e-19
C12 clk gnd 0.030199f
C13 qbar clk 6.44e-19
C14 vdd a_n206_n60# 0.41238f
C15 w_n216_n73# a_n214_n85# 0.04795f
C16 a_n137_n36# gnd 7.27e-19
C17 a_n214_n85# gnd 0.20619f
C18 d clk 0.041238f
C19 vdd a_n137_n36# 0.41238f
C20 w_n216_n43# vdd 0.008089f
C21 a_n144_n85# gnd 0.20619f
C22 a_n206_n60# clk 0.020744f
C23 w_n147_n43# vdd 0.006878f
C24 w_n216_n43# d 0.026794f
C25 w_n85_n43# qbar 0.007278f
C26 a_n82_n85# gnd 0.20619f
C27 w_n23_n70# q 0.013119f
C28 qbar a_n82_n85# 0.318127f
C29 w_n216_n43# a_n206_n60# 0.007029f
C30 w_n85_n43# vdd 0.006926f
C31 q gnd 0.20619f
C32 a_n206_n60# a_n214_n85# 0.453629f
C33 clk a_n137_n36# 0.013701f
C34 qbar q 0.062736f
C35 w_n23_n70# qbar 0.027447f
C36 w_n216_n43# clk 4.5e-19
C37 qbar gnd 0.042287f
C38 vdd q 0.439883f
C39 clk a_n214_n85# 0.033079f
C40 w_n147_n43# clk 0.027431f
C41 w_n23_n70# vdd 0.008693f
C42 gnd 0 0.796845f  
C43 q 0 0.165505f  
C44 a_n82_n85# 0 0.170919f  
C45 a_n144_n85# 0 0.20023f  
C46 a_n214_n85# 0 0.356257f  
C47 a_n137_n36# 0 0.476334f  
C48 clk 0 3.22455f  
C49 a_n206_n60# 0 0.128632f  
C50 d 0 0.470088f  
C51 vdd 0 0.77082f  
C52 qbar 0 0.51689f  
C53 w_n23_n70# 0 1.68739f  
C54 w_n216_n73# 0 1.34991f  
C55 w_n85_n43# 0 1.40616f  
C56 w_n147_n43# 0 1.40616f  
C57 w_n216_n43# 0 1.40616f  






.control
  set hcopypscolor = 1
  set color0 = white
  set color1 = black
  set color2 = red
  set color3 = blue
  set color4 = green
  set color5 = brown
  set color6 = magenta
  set color7 = cyan
  tran 1n 200n
  plot clk d+2 q+4 qbar+6 
  * Measure propagation delay from D to Q_actual
  meas tran tpd_d_q_actual_rise TRIG v(d) VAL=0.9 RISE=1 TARG v(q) VAL=0.9 RISE=1
  meas tran tpd_d_q_actual_fall TRIG v(d) VAL=0.9 FALL=1 TARG v(q) VAL=0.9 FALL=1
  let delay_d_q_actual = abs((tpd_d_q_actual_rise + tpd_d_q_actual_fall)/2)
  print delay_d_q_actual

  * Measure rise and fall times of Q_actual
  meas tran tr_q_actual TRIG v(q) VAL=0.9 RISE=1 TARG v(q) VAL=1.8 RISE=1
  meas tran tf_q_actual TRIG v(q) VAL=1.8 FALL=1 TARG v(q) VAL=0.9 FALL=1
  print tr_q_actual tf_q_actual

  * Measure setup and hold times
  meas tran t_setup TRIG v(clk) VAL=0.9 RISE=1 TARG v(d) VAL=0.9 FALL=1
  meas tran t_hold TRIG v(clk) VAL=0.9 RISE=1 TARG v(d) VAL=0.9 RISE=1
  print t_setup t_hold
.endc
.end
