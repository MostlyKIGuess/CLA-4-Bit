magic
tech scmos
timestamp 1731837759
<< nwell >>
rect 193 588 217 644
rect 226 594 250 650
rect 302 599 326 655
rect 335 599 359 655
rect 368 604 392 660
rect 401 604 425 660
rect 434 604 458 660
rect 472 604 496 660
rect 505 625 529 681
rect 538 625 562 681
rect 571 625 595 681
rect 604 625 628 681
rect 642 625 666 681
rect 675 654 699 710
rect 708 654 732 710
rect 741 654 765 710
rect 774 654 798 710
rect 807 654 831 710
rect 845 654 869 710
rect 205 450 229 506
rect 238 456 262 512
rect 314 461 338 517
rect 347 461 371 517
rect 384 462 408 518
rect 417 462 441 518
rect 450 462 474 518
rect 488 462 512 518
rect 521 464 545 520
rect 554 464 578 520
rect 587 464 611 520
rect 620 464 644 520
rect 658 464 682 520
rect 726 513 782 537
rect 879 518 935 542
rect 725 479 781 503
rect 878 485 934 509
rect 725 444 781 468
rect -108 412 -52 437
rect -39 412 17 437
rect 23 412 79 437
rect -108 382 -52 406
rect 85 385 115 441
rect 725 411 781 435
rect 790 410 814 466
rect 877 451 933 475
rect 1035 443 1091 468
rect 1104 443 1160 468
rect 1166 443 1222 468
rect 877 416 933 440
rect 877 383 933 407
rect 942 382 966 438
rect 1035 413 1091 437
rect 1228 416 1258 472
rect -109 298 -53 323
rect -40 298 16 323
rect 22 298 78 323
rect -109 268 -53 292
rect 84 271 114 327
rect 258 312 282 368
rect 291 318 315 374
rect 367 323 391 379
rect 400 323 424 379
rect 440 301 464 357
rect 473 301 497 357
rect 506 301 530 357
rect 544 301 568 357
rect 611 340 667 364
rect 611 305 667 329
rect 611 272 667 296
rect 676 271 700 327
rect 725 266 749 322
rect 758 272 782 328
rect 797 280 821 332
rect 834 277 858 333
rect 867 277 891 333
rect -106 184 -50 209
rect -37 184 19 209
rect 25 184 81 209
rect -106 154 -50 178
rect 87 157 117 213
rect 258 174 282 230
rect 291 180 315 236
rect 367 185 391 241
rect 400 185 424 241
rect 439 167 495 191
rect 439 134 495 158
rect 504 133 528 189
rect -103 70 -47 95
rect -34 70 22 95
rect 28 70 84 95
rect -103 40 -47 64
rect 90 43 120 99
rect 258 17 282 73
rect 291 17 315 73
rect 328 18 352 70
rect 367 22 391 78
rect 400 28 424 84
rect 551 57 575 113
rect 584 63 608 119
rect 660 68 684 124
rect 693 68 717 124
rect 1016 123 1072 148
rect 1085 123 1141 148
rect 1147 123 1203 148
rect 1016 93 1072 117
rect 1209 96 1239 152
rect 1015 9 1071 34
rect 1084 9 1140 34
rect 1146 9 1202 34
rect -104 -48 -48 -23
rect -35 -48 21 -23
rect 27 -48 83 -23
rect -104 -78 -48 -54
rect 89 -75 119 -19
rect 258 -117 282 -61
rect 291 -117 315 -61
rect 328 -116 352 -64
rect 367 -112 391 -56
rect 400 -106 424 -50
rect 548 -81 572 -25
rect 581 -75 605 -19
rect 657 -70 681 -14
rect 690 -70 714 -14
rect 785 -81 809 -25
rect 818 -75 842 -19
rect 857 -67 881 -15
rect 1015 -21 1071 3
rect 1208 -18 1238 38
rect 1018 -105 1074 -80
rect 1087 -105 1143 -80
rect 1149 -105 1205 -80
rect -105 -162 -49 -137
rect -36 -162 20 -137
rect 26 -162 82 -137
rect -105 -192 -49 -168
rect 88 -189 118 -133
rect 1018 -135 1074 -111
rect 1211 -132 1241 -76
rect -102 -276 -46 -251
rect -33 -276 23 -251
rect 29 -276 85 -251
rect -102 -306 -46 -282
rect 91 -303 121 -247
rect 329 -250 353 -198
rect 368 -246 392 -190
rect 401 -240 425 -184
rect 551 -219 575 -163
rect 584 -213 608 -157
rect 782 -215 806 -159
rect 815 -209 839 -153
rect 854 -201 878 -149
rect 1021 -219 1077 -194
rect 1090 -219 1146 -194
rect 1152 -219 1208 -194
rect 1021 -249 1077 -225
rect 1214 -246 1244 -190
rect -99 -390 -43 -365
rect -30 -390 26 -365
rect 32 -390 88 -365
rect -99 -420 -43 -396
rect 94 -417 124 -361
rect 329 -384 353 -332
rect 368 -380 392 -324
rect 401 -374 425 -318
rect 551 -357 575 -301
rect 584 -351 608 -295
rect 660 -346 684 -290
rect 693 -346 717 -290
rect 795 -349 819 -293
rect 828 -343 852 -287
rect 867 -335 891 -283
<< ntransistor >>
rect 252 667 272 669
rect 797 621 837 623
rect 856 622 858 642
rect 252 581 272 583
rect 204 556 206 576
rect 313 567 315 587
rect 346 567 348 587
rect 424 571 464 573
rect 483 572 485 592
rect 594 592 634 594
rect 653 593 655 613
rect 797 602 837 604
rect 797 583 837 585
rect 594 573 634 575
rect 797 564 837 566
rect 424 552 464 554
rect 594 554 634 556
rect 797 545 837 547
rect 424 533 464 535
rect 594 535 634 537
rect 264 529 284 531
rect 264 443 284 445
rect -10 399 10 401
rect 52 399 72 401
rect 216 418 218 438
rect 325 429 327 449
rect 358 429 360 449
rect 440 429 480 431
rect 499 430 501 450
rect 610 431 650 433
rect 669 432 671 452
rect 440 410 480 412
rect 610 412 650 414
rect -106 368 -86 370
rect -36 368 -16 370
rect 26 368 46 370
rect 317 391 337 393
rect 440 391 480 393
rect 610 393 650 395
rect 691 378 693 398
rect 712 378 714 398
rect 741 378 743 398
rect 774 378 776 398
rect 801 378 803 398
rect 1133 430 1153 432
rect 1195 430 1215 432
rect 1037 399 1057 401
rect 1107 399 1127 401
rect 1169 399 1189 401
rect 610 375 650 377
rect 102 345 104 365
rect 1245 376 1247 396
rect -11 285 9 287
rect 51 285 71 287
rect 823 350 825 370
rect 843 350 845 370
rect 864 350 866 370
rect 893 350 895 370
rect 926 350 928 370
rect 953 350 955 370
rect 317 305 337 307
rect -107 254 -87 256
rect -37 254 -17 256
rect 25 254 45 256
rect 269 280 271 300
rect 378 291 380 311
rect 411 291 413 311
rect 496 268 536 270
rect 555 269 557 289
rect 317 253 337 255
rect 101 231 103 251
rect 496 249 536 251
rect 598 239 600 259
rect 627 239 629 259
rect 660 239 662 259
rect 687 239 689 259
rect 784 258 804 260
rect -8 171 12 173
rect 54 171 74 173
rect 736 234 738 254
rect 496 230 536 232
rect 821 233 823 253
rect 845 245 847 265
rect 878 245 880 265
rect -104 140 -84 142
rect -34 140 -14 142
rect 28 140 48 142
rect 317 167 337 169
rect 269 142 271 162
rect 378 153 380 173
rect 411 153 413 173
rect 104 117 106 137
rect 610 136 630 138
rect -5 57 15 59
rect 57 57 77 59
rect 269 85 271 105
rect 302 85 304 105
rect 326 97 328 117
rect 411 96 413 116
rect 455 101 457 121
rect 488 101 490 121
rect 515 101 517 121
rect 345 90 365 92
rect -101 26 -81 28
rect -31 26 -11 28
rect 31 26 51 28
rect 1114 110 1134 112
rect 1176 110 1196 112
rect 1018 79 1038 81
rect 1088 79 1108 81
rect 1150 79 1170 81
rect 1226 56 1228 76
rect 610 50 630 52
rect 562 25 564 45
rect 671 36 673 56
rect 704 36 706 56
rect 107 3 109 23
rect 607 -2 627 0
rect 1113 -4 1133 -2
rect 1175 -4 1195 -2
rect -6 -61 14 -59
rect 56 -61 76 -59
rect 269 -49 271 -29
rect 302 -49 304 -29
rect 326 -37 328 -17
rect 411 -38 413 -18
rect 345 -44 365 -42
rect -102 -92 -82 -90
rect -32 -92 -12 -90
rect 30 -92 50 -90
rect 106 -115 108 -95
rect 1017 -35 1037 -33
rect 1087 -35 1107 -33
rect 1149 -35 1169 -33
rect 1225 -58 1227 -38
rect 607 -88 627 -86
rect 559 -113 561 -93
rect 668 -102 670 -82
rect 701 -102 703 -82
rect 844 -89 864 -87
rect 796 -113 798 -93
rect 881 -114 883 -94
rect 1116 -118 1136 -116
rect 1178 -118 1198 -116
rect -7 -175 13 -173
rect 55 -175 75 -173
rect 610 -140 630 -138
rect 327 -171 329 -151
rect 1020 -149 1040 -147
rect 1090 -149 1110 -147
rect 1152 -149 1172 -147
rect 412 -172 414 -152
rect -103 -206 -83 -204
rect -33 -206 -13 -204
rect 29 -206 49 -204
rect 346 -178 366 -176
rect 105 -229 107 -209
rect 1228 -172 1230 -152
rect 610 -226 630 -224
rect 841 -223 861 -221
rect 562 -251 564 -231
rect 793 -247 795 -227
rect 878 -248 880 -228
rect 1119 -232 1139 -230
rect 1181 -232 1201 -230
rect -4 -289 16 -287
rect 58 -289 78 -287
rect 1023 -263 1043 -261
rect 1093 -263 1113 -261
rect 1155 -263 1175 -261
rect 610 -278 630 -276
rect -100 -320 -80 -318
rect -30 -320 -10 -318
rect 32 -320 52 -318
rect 327 -305 329 -285
rect 1231 -286 1233 -266
rect 412 -306 414 -286
rect 346 -312 366 -310
rect 108 -343 110 -323
rect -1 -403 19 -401
rect 61 -403 81 -401
rect 610 -364 630 -362
rect 562 -389 564 -369
rect 671 -378 673 -358
rect 704 -378 706 -358
rect 854 -357 874 -355
rect 806 -381 808 -361
rect 891 -382 893 -362
rect -97 -434 -77 -432
rect -27 -434 -7 -432
rect 35 -434 55 -432
rect 111 -457 113 -437
<< ptransistor >>
rect 204 598 206 638
rect 237 604 239 644
rect 313 609 315 649
rect 346 609 348 649
rect 379 614 381 654
rect 412 614 414 654
rect 445 614 447 654
rect 483 614 485 654
rect 516 635 518 675
rect 549 635 551 675
rect 582 635 584 675
rect 615 635 617 675
rect 653 635 655 675
rect 686 664 688 704
rect 719 664 721 704
rect 752 664 754 704
rect 785 664 787 704
rect 818 664 820 704
rect 856 664 858 704
rect 885 529 925 531
rect 732 524 772 526
rect 216 460 218 500
rect 249 466 251 506
rect 325 471 327 511
rect 358 471 360 511
rect 395 472 397 512
rect 428 472 430 512
rect 461 472 463 512
rect 499 472 501 512
rect 532 474 534 514
rect 565 474 567 514
rect 598 474 600 514
rect 631 474 633 514
rect 669 474 671 514
rect 884 496 924 498
rect 731 490 771 492
rect 883 462 923 464
rect 731 455 771 457
rect -98 424 -58 426
rect -29 424 11 426
rect 33 424 73 426
rect -98 393 -58 395
rect 102 395 104 435
rect 731 422 771 424
rect 801 420 803 460
rect 1045 455 1085 457
rect 1114 455 1154 457
rect 1176 455 1216 457
rect 883 427 923 429
rect 883 394 923 396
rect 953 392 955 432
rect 1045 424 1085 426
rect 1245 426 1247 466
rect 269 322 271 362
rect 302 328 304 368
rect 378 333 380 373
rect 411 333 413 373
rect -99 310 -59 312
rect -30 310 10 312
rect 32 310 72 312
rect -99 279 -59 281
rect 101 281 103 321
rect 451 311 453 351
rect 484 311 486 351
rect 517 311 519 351
rect 555 311 557 351
rect 617 351 657 353
rect 617 316 657 318
rect 617 283 657 285
rect 687 281 689 321
rect 736 276 738 316
rect 769 282 771 322
rect 808 286 810 326
rect 845 287 847 327
rect 878 287 880 327
rect -96 196 -56 198
rect -27 196 13 198
rect 35 196 75 198
rect -96 165 -56 167
rect 104 167 106 207
rect 269 184 271 224
rect 302 190 304 230
rect 378 195 380 235
rect 411 195 413 235
rect 445 178 485 180
rect 445 145 485 147
rect 515 143 517 183
rect 1026 135 1066 137
rect 1095 135 1135 137
rect 1157 135 1197 137
rect -93 82 -53 84
rect -24 82 16 84
rect 38 82 78 84
rect -93 51 -53 53
rect 107 53 109 93
rect 269 23 271 63
rect 302 23 304 63
rect 339 24 341 64
rect 378 28 380 68
rect 411 34 413 74
rect 562 67 564 107
rect 595 73 597 113
rect 671 78 673 118
rect 704 78 706 118
rect 1026 104 1066 106
rect 1226 106 1228 146
rect 1025 21 1065 23
rect 1094 21 1134 23
rect 1156 21 1196 23
rect 1025 -10 1065 -8
rect 1225 -8 1227 32
rect -94 -36 -54 -34
rect -25 -36 15 -34
rect 37 -36 77 -34
rect -94 -67 -54 -65
rect 106 -65 108 -25
rect 269 -111 271 -71
rect 302 -111 304 -71
rect 339 -110 341 -70
rect 378 -106 380 -66
rect 411 -100 413 -60
rect 559 -71 561 -31
rect 592 -65 594 -25
rect 668 -60 670 -20
rect 701 -60 703 -20
rect 796 -71 798 -31
rect 829 -65 831 -25
rect 868 -61 870 -21
rect 1028 -93 1068 -91
rect 1097 -93 1137 -91
rect 1159 -93 1199 -91
rect 1028 -124 1068 -122
rect 1228 -122 1230 -82
rect -95 -150 -55 -148
rect -26 -150 14 -148
rect 36 -150 76 -148
rect -95 -181 -55 -179
rect 105 -179 107 -139
rect 340 -244 342 -204
rect 379 -240 381 -200
rect 412 -234 414 -194
rect 562 -209 564 -169
rect 595 -203 597 -163
rect 793 -205 795 -165
rect 826 -199 828 -159
rect 865 -195 867 -155
rect 1031 -207 1071 -205
rect 1100 -207 1140 -205
rect 1162 -207 1202 -205
rect 1031 -238 1071 -236
rect 1231 -236 1233 -196
rect -92 -264 -52 -262
rect -23 -264 17 -262
rect 39 -264 79 -262
rect -92 -295 -52 -293
rect 108 -293 110 -253
rect -89 -378 -49 -376
rect -20 -378 20 -376
rect 42 -378 82 -376
rect -89 -409 -49 -407
rect 111 -407 113 -367
rect 340 -378 342 -338
rect 379 -374 381 -334
rect 412 -368 414 -328
rect 562 -347 564 -307
rect 595 -341 597 -301
rect 671 -336 673 -296
rect 704 -336 706 -296
rect 806 -339 808 -299
rect 839 -333 841 -293
rect 878 -329 880 -289
<< ndiffusion >>
rect 252 669 272 670
rect 252 666 272 667
rect 797 623 837 624
rect 855 622 856 642
rect 858 622 859 642
rect 797 620 837 621
rect 252 583 272 584
rect 252 580 272 581
rect 203 556 204 576
rect 206 556 207 576
rect 312 567 313 587
rect 315 567 316 587
rect 345 567 346 587
rect 348 567 349 587
rect 424 573 464 574
rect 482 572 483 592
rect 485 572 486 592
rect 594 594 634 595
rect 652 593 653 613
rect 655 593 656 613
rect 797 604 837 605
rect 797 601 837 602
rect 594 591 634 592
rect 797 585 837 586
rect 797 582 837 583
rect 424 570 464 571
rect 594 575 634 576
rect 594 572 634 573
rect 797 566 837 567
rect 797 563 837 564
rect 424 554 464 555
rect 594 556 634 557
rect 594 553 634 554
rect 424 551 464 552
rect 797 547 837 548
rect 797 544 837 545
rect 264 531 284 532
rect 424 535 464 536
rect 594 537 634 538
rect 594 534 634 535
rect 424 532 464 533
rect 264 528 284 529
rect 264 445 284 446
rect 264 442 284 443
rect -10 401 10 402
rect -10 398 10 399
rect 52 401 72 402
rect 52 398 72 399
rect 215 418 216 438
rect 218 418 219 438
rect 324 429 325 449
rect 327 429 328 449
rect 357 429 358 449
rect 360 429 361 449
rect 440 431 480 432
rect 498 430 499 450
rect 501 430 502 450
rect 440 428 480 429
rect 610 433 650 434
rect 668 432 669 452
rect 671 432 672 452
rect 610 430 650 431
rect 440 412 480 413
rect 610 414 650 415
rect 610 411 650 412
rect 440 409 480 410
rect -106 370 -86 371
rect -106 367 -86 368
rect -36 370 -16 371
rect 26 370 46 371
rect -36 367 -16 368
rect 26 367 46 368
rect 317 393 337 394
rect 317 390 337 391
rect 440 393 480 394
rect 610 395 650 396
rect 610 392 650 393
rect 440 390 480 391
rect 690 378 691 398
rect 693 378 694 398
rect 711 378 712 398
rect 714 378 715 398
rect 740 378 741 398
rect 743 378 744 398
rect 773 378 774 398
rect 776 378 777 398
rect 800 378 801 398
rect 803 378 804 398
rect 1133 432 1153 433
rect 1133 429 1153 430
rect 1195 432 1215 433
rect 1195 429 1215 430
rect 1037 401 1057 402
rect 1037 398 1057 399
rect 1107 401 1127 402
rect 1169 401 1189 402
rect 1107 398 1127 399
rect 1169 398 1189 399
rect 610 377 650 378
rect 610 374 650 375
rect 101 345 102 365
rect 104 345 105 365
rect 1244 376 1245 396
rect 1247 376 1248 396
rect -11 287 9 288
rect -11 284 9 285
rect 51 287 71 288
rect 51 284 71 285
rect 822 350 823 370
rect 825 350 826 370
rect 842 350 843 370
rect 845 350 846 370
rect 863 350 864 370
rect 866 350 867 370
rect 892 350 893 370
rect 895 350 896 370
rect 925 350 926 370
rect 928 350 929 370
rect 952 350 953 370
rect 955 350 956 370
rect 317 307 337 308
rect 317 304 337 305
rect -107 256 -87 257
rect -107 253 -87 254
rect -37 256 -17 257
rect 25 256 45 257
rect -37 253 -17 254
rect 25 253 45 254
rect 268 280 269 300
rect 271 280 272 300
rect 377 291 378 311
rect 380 291 381 311
rect 410 291 411 311
rect 413 291 414 311
rect 496 270 536 271
rect 554 269 555 289
rect 557 269 558 289
rect 496 267 536 268
rect 317 255 337 256
rect 317 252 337 253
rect 100 231 101 251
rect 103 231 104 251
rect 496 251 536 252
rect 496 248 536 249
rect 597 239 598 259
rect 600 239 601 259
rect 626 239 627 259
rect 629 239 630 259
rect 659 239 660 259
rect 662 239 663 259
rect 686 239 687 259
rect 689 239 690 259
rect 784 260 804 261
rect 784 257 804 258
rect -8 173 12 174
rect -8 170 12 171
rect 54 173 74 174
rect 54 170 74 171
rect 735 234 736 254
rect 738 234 739 254
rect 496 232 536 233
rect 820 233 821 253
rect 823 233 824 253
rect 844 245 845 265
rect 847 245 848 265
rect 877 245 878 265
rect 880 245 881 265
rect 496 229 536 230
rect -104 142 -84 143
rect -104 139 -84 140
rect -34 142 -14 143
rect 28 142 48 143
rect -34 139 -14 140
rect 28 139 48 140
rect 317 169 337 170
rect 317 166 337 167
rect 268 142 269 162
rect 271 142 272 162
rect 377 153 378 173
rect 380 153 381 173
rect 410 153 411 173
rect 413 153 414 173
rect 103 117 104 137
rect 106 117 107 137
rect 610 138 630 139
rect 610 135 630 136
rect -5 59 15 60
rect -5 56 15 57
rect 57 59 77 60
rect 57 56 77 57
rect 268 85 269 105
rect 271 85 272 105
rect 301 85 302 105
rect 304 85 305 105
rect 325 97 326 117
rect 328 97 329 117
rect 410 96 411 116
rect 413 96 414 116
rect 454 101 455 121
rect 457 101 458 121
rect 487 101 488 121
rect 490 101 491 121
rect 514 101 515 121
rect 517 101 518 121
rect 345 92 365 93
rect 345 89 365 90
rect -101 28 -81 29
rect -101 25 -81 26
rect -31 28 -11 29
rect 31 28 51 29
rect -31 25 -11 26
rect 31 25 51 26
rect 1114 112 1134 113
rect 1114 109 1134 110
rect 1176 112 1196 113
rect 1176 109 1196 110
rect 1018 81 1038 82
rect 1018 78 1038 79
rect 1088 81 1108 82
rect 1150 81 1170 82
rect 1088 78 1108 79
rect 1150 78 1170 79
rect 1225 56 1226 76
rect 1228 56 1229 76
rect 610 52 630 53
rect 610 49 630 50
rect 561 25 562 45
rect 564 25 565 45
rect 670 36 671 56
rect 673 36 674 56
rect 703 36 704 56
rect 706 36 707 56
rect 106 3 107 23
rect 109 3 110 23
rect 607 0 627 1
rect 607 -3 627 -2
rect 1113 -2 1133 -1
rect 1113 -5 1133 -4
rect 1175 -2 1195 -1
rect 1175 -5 1195 -4
rect -6 -59 14 -58
rect -6 -62 14 -61
rect 56 -59 76 -58
rect 56 -62 76 -61
rect 268 -49 269 -29
rect 271 -49 272 -29
rect 301 -49 302 -29
rect 304 -49 305 -29
rect 325 -37 326 -17
rect 328 -37 329 -17
rect 410 -38 411 -18
rect 413 -38 414 -18
rect 345 -42 365 -41
rect 345 -45 365 -44
rect -102 -90 -82 -89
rect -102 -93 -82 -92
rect -32 -90 -12 -89
rect 30 -90 50 -89
rect -32 -93 -12 -92
rect 30 -93 50 -92
rect 105 -115 106 -95
rect 108 -115 109 -95
rect 1017 -33 1037 -32
rect 1017 -36 1037 -35
rect 1087 -33 1107 -32
rect 1149 -33 1169 -32
rect 1087 -36 1107 -35
rect 1149 -36 1169 -35
rect 1224 -58 1225 -38
rect 1227 -58 1228 -38
rect 607 -86 627 -85
rect 607 -89 627 -88
rect 558 -113 559 -93
rect 561 -113 562 -93
rect 667 -102 668 -82
rect 670 -102 671 -82
rect 700 -102 701 -82
rect 703 -102 704 -82
rect 844 -87 864 -86
rect 844 -90 864 -89
rect 795 -113 796 -93
rect 798 -113 799 -93
rect 880 -114 881 -94
rect 883 -114 884 -94
rect 1116 -116 1136 -115
rect 1116 -119 1136 -118
rect 1178 -116 1198 -115
rect 1178 -119 1198 -118
rect -7 -173 13 -172
rect -7 -176 13 -175
rect 55 -173 75 -172
rect 55 -176 75 -175
rect 610 -138 630 -137
rect 610 -141 630 -140
rect 326 -171 327 -151
rect 329 -171 330 -151
rect 1020 -147 1040 -146
rect 1020 -150 1040 -149
rect 1090 -147 1110 -146
rect 1152 -147 1172 -146
rect 1090 -150 1110 -149
rect 411 -172 412 -152
rect 414 -172 415 -152
rect 1152 -150 1172 -149
rect -103 -204 -83 -203
rect -103 -207 -83 -206
rect -33 -204 -13 -203
rect 29 -204 49 -203
rect -33 -207 -13 -206
rect 29 -207 49 -206
rect 346 -176 366 -175
rect 346 -179 366 -178
rect 104 -229 105 -209
rect 107 -229 108 -209
rect 1227 -172 1228 -152
rect 1230 -172 1231 -152
rect 610 -224 630 -223
rect 610 -227 630 -226
rect 841 -221 861 -220
rect 841 -224 861 -223
rect 561 -251 562 -231
rect 564 -251 565 -231
rect 792 -247 793 -227
rect 795 -247 796 -227
rect 877 -248 878 -228
rect 880 -248 881 -228
rect 1119 -230 1139 -229
rect 1119 -233 1139 -232
rect 1181 -230 1201 -229
rect 1181 -233 1201 -232
rect -4 -287 16 -286
rect -4 -290 16 -289
rect 58 -287 78 -286
rect 58 -290 78 -289
rect 1023 -261 1043 -260
rect 1023 -264 1043 -263
rect 1093 -261 1113 -260
rect 1155 -261 1175 -260
rect 1093 -264 1113 -263
rect 1155 -264 1175 -263
rect 610 -276 630 -275
rect 610 -279 630 -278
rect -100 -318 -80 -317
rect -100 -321 -80 -320
rect -30 -318 -10 -317
rect 32 -318 52 -317
rect -30 -321 -10 -320
rect 32 -321 52 -320
rect 326 -305 327 -285
rect 329 -305 330 -285
rect 1230 -286 1231 -266
rect 1233 -286 1234 -266
rect 411 -306 412 -286
rect 414 -306 415 -286
rect 346 -310 366 -309
rect 346 -313 366 -312
rect 107 -343 108 -323
rect 110 -343 111 -323
rect -1 -401 19 -400
rect -1 -404 19 -403
rect 61 -401 81 -400
rect 61 -404 81 -403
rect 610 -362 630 -361
rect 610 -365 630 -364
rect 561 -389 562 -369
rect 564 -389 565 -369
rect 670 -378 671 -358
rect 673 -378 674 -358
rect 703 -378 704 -358
rect 706 -378 707 -358
rect 854 -355 874 -354
rect 854 -358 874 -357
rect 805 -381 806 -361
rect 808 -381 809 -361
rect 890 -382 891 -362
rect 893 -382 894 -362
rect -97 -432 -77 -431
rect -97 -435 -77 -434
rect -27 -432 -7 -431
rect 35 -432 55 -431
rect -27 -435 -7 -434
rect 35 -435 55 -434
rect 110 -457 111 -437
rect 113 -457 114 -437
<< pdiffusion >>
rect 203 598 204 638
rect 206 598 207 638
rect 236 604 237 644
rect 239 604 240 644
rect 312 609 313 649
rect 315 609 316 649
rect 345 609 346 649
rect 348 609 349 649
rect 378 614 379 654
rect 381 614 382 654
rect 411 614 412 654
rect 414 614 415 654
rect 444 614 445 654
rect 447 614 448 654
rect 482 614 483 654
rect 485 614 486 654
rect 515 635 516 675
rect 518 635 519 675
rect 548 635 549 675
rect 551 635 552 675
rect 581 635 582 675
rect 584 635 585 675
rect 614 635 615 675
rect 617 635 618 675
rect 652 635 653 675
rect 655 635 656 675
rect 685 664 686 704
rect 688 664 689 704
rect 718 664 719 704
rect 721 664 722 704
rect 751 664 752 704
rect 754 664 755 704
rect 784 664 785 704
rect 787 664 788 704
rect 817 664 818 704
rect 820 664 821 704
rect 855 664 856 704
rect 858 664 859 704
rect 885 531 925 532
rect 885 528 925 529
rect 732 526 772 527
rect 732 523 772 524
rect 215 460 216 500
rect 218 460 219 500
rect 248 466 249 506
rect 251 466 252 506
rect 324 471 325 511
rect 327 471 328 511
rect 357 471 358 511
rect 360 471 361 511
rect 394 472 395 512
rect 397 472 398 512
rect 427 472 428 512
rect 430 472 431 512
rect 460 472 461 512
rect 463 472 464 512
rect 498 472 499 512
rect 501 472 502 512
rect 531 474 532 514
rect 534 474 535 514
rect 564 474 565 514
rect 567 474 568 514
rect 597 474 598 514
rect 600 474 601 514
rect 630 474 631 514
rect 633 474 634 514
rect 668 474 669 514
rect 671 474 672 514
rect 884 498 924 499
rect 884 495 924 496
rect 731 492 771 493
rect 731 489 771 490
rect 883 464 923 465
rect 883 461 923 462
rect 731 457 771 458
rect 731 454 771 455
rect -98 426 -58 427
rect -98 423 -58 424
rect -29 426 11 427
rect -29 423 11 424
rect 33 426 73 427
rect 33 423 73 424
rect -98 395 -58 396
rect 101 395 102 435
rect 104 395 105 435
rect 731 424 771 425
rect 731 421 771 422
rect 800 420 801 460
rect 803 420 804 460
rect 1045 457 1085 458
rect 1045 454 1085 455
rect 1114 457 1154 458
rect 1114 454 1154 455
rect 1176 457 1216 458
rect 1176 454 1216 455
rect 883 429 923 430
rect 883 426 923 427
rect -98 392 -58 393
rect 883 396 923 397
rect 883 393 923 394
rect 952 392 953 432
rect 955 392 956 432
rect 1045 426 1085 427
rect 1244 426 1245 466
rect 1247 426 1248 466
rect 1045 423 1085 424
rect 268 322 269 362
rect 271 322 272 362
rect 301 328 302 368
rect 304 328 305 368
rect 377 333 378 373
rect 380 333 381 373
rect 410 333 411 373
rect 413 333 414 373
rect -99 312 -59 313
rect -99 309 -59 310
rect -30 312 10 313
rect -30 309 10 310
rect 32 312 72 313
rect 32 309 72 310
rect -99 281 -59 282
rect 100 281 101 321
rect 103 281 104 321
rect 450 311 451 351
rect 453 311 454 351
rect 483 311 484 351
rect 486 311 487 351
rect 516 311 517 351
rect 519 311 520 351
rect 554 311 555 351
rect 557 311 558 351
rect 617 353 657 354
rect 617 350 657 351
rect 617 318 657 319
rect 617 315 657 316
rect -99 278 -59 279
rect 617 285 657 286
rect 617 282 657 283
rect 686 281 687 321
rect 689 281 690 321
rect 735 276 736 316
rect 738 276 739 316
rect 768 282 769 322
rect 771 282 772 322
rect 807 286 808 326
rect 810 286 811 326
rect 844 287 845 327
rect 847 287 848 327
rect 877 287 878 327
rect 880 287 881 327
rect -96 198 -56 199
rect -96 195 -56 196
rect -27 198 13 199
rect -27 195 13 196
rect 35 198 75 199
rect 35 195 75 196
rect -96 167 -56 168
rect 103 167 104 207
rect 106 167 107 207
rect 268 184 269 224
rect 271 184 272 224
rect 301 190 302 230
rect 304 190 305 230
rect 377 195 378 235
rect 380 195 381 235
rect 410 195 411 235
rect 413 195 414 235
rect -96 164 -56 165
rect 445 180 485 181
rect 445 177 485 178
rect 445 147 485 148
rect 445 144 485 145
rect 514 143 515 183
rect 517 143 518 183
rect 1026 137 1066 138
rect 1026 134 1066 135
rect 1095 137 1135 138
rect 1095 134 1135 135
rect 1157 137 1197 138
rect 1157 134 1197 135
rect -93 84 -53 85
rect -93 81 -53 82
rect -24 84 16 85
rect -24 81 16 82
rect 38 84 78 85
rect 38 81 78 82
rect -93 53 -53 54
rect 106 53 107 93
rect 109 53 110 93
rect -93 50 -53 51
rect 268 23 269 63
rect 271 23 272 63
rect 301 23 302 63
rect 304 23 305 63
rect 338 24 339 64
rect 341 24 342 64
rect 377 28 378 68
rect 380 28 381 68
rect 410 34 411 74
rect 413 34 414 74
rect 561 67 562 107
rect 564 67 565 107
rect 594 73 595 113
rect 597 73 598 113
rect 670 78 671 118
rect 673 78 674 118
rect 703 78 704 118
rect 706 78 707 118
rect 1026 106 1066 107
rect 1225 106 1226 146
rect 1228 106 1229 146
rect 1026 103 1066 104
rect 1025 23 1065 24
rect 1025 20 1065 21
rect 1094 23 1134 24
rect 1094 20 1134 21
rect 1156 23 1196 24
rect 1156 20 1196 21
rect 1025 -8 1065 -7
rect 1224 -8 1225 32
rect 1227 -8 1228 32
rect 1025 -11 1065 -10
rect -94 -34 -54 -33
rect -94 -37 -54 -36
rect -25 -34 15 -33
rect -25 -37 15 -36
rect 37 -34 77 -33
rect 37 -37 77 -36
rect -94 -65 -54 -64
rect 105 -65 106 -25
rect 108 -65 109 -25
rect -94 -68 -54 -67
rect 268 -111 269 -71
rect 271 -111 272 -71
rect 301 -111 302 -71
rect 304 -111 305 -71
rect 338 -110 339 -70
rect 341 -110 342 -70
rect 377 -106 378 -66
rect 380 -106 381 -66
rect 410 -100 411 -60
rect 413 -100 414 -60
rect 558 -71 559 -31
rect 561 -71 562 -31
rect 591 -65 592 -25
rect 594 -65 595 -25
rect 667 -60 668 -20
rect 670 -60 671 -20
rect 700 -60 701 -20
rect 703 -60 704 -20
rect 795 -71 796 -31
rect 798 -71 799 -31
rect 828 -65 829 -25
rect 831 -65 832 -25
rect 867 -61 868 -21
rect 870 -61 871 -21
rect 1028 -91 1068 -90
rect 1028 -94 1068 -93
rect 1097 -91 1137 -90
rect 1097 -94 1137 -93
rect 1159 -91 1199 -90
rect 1159 -94 1199 -93
rect 1028 -122 1068 -121
rect 1227 -122 1228 -82
rect 1230 -122 1231 -82
rect 1028 -125 1068 -124
rect -95 -148 -55 -147
rect -95 -151 -55 -150
rect -26 -148 14 -147
rect -26 -151 14 -150
rect 36 -148 76 -147
rect 36 -151 76 -150
rect -95 -179 -55 -178
rect 104 -179 105 -139
rect 107 -179 108 -139
rect -95 -182 -55 -181
rect 339 -244 340 -204
rect 342 -244 343 -204
rect 378 -240 379 -200
rect 381 -240 382 -200
rect 411 -234 412 -194
rect 414 -234 415 -194
rect 561 -209 562 -169
rect 564 -209 565 -169
rect 594 -203 595 -163
rect 597 -203 598 -163
rect 792 -205 793 -165
rect 795 -205 796 -165
rect 825 -199 826 -159
rect 828 -199 829 -159
rect 864 -195 865 -155
rect 867 -195 868 -155
rect 1031 -205 1071 -204
rect 1031 -208 1071 -207
rect 1100 -205 1140 -204
rect 1100 -208 1140 -207
rect 1162 -205 1202 -204
rect 1162 -208 1202 -207
rect 1031 -236 1071 -235
rect 1230 -236 1231 -196
rect 1233 -236 1234 -196
rect 1031 -239 1071 -238
rect -92 -262 -52 -261
rect -92 -265 -52 -264
rect -23 -262 17 -261
rect -23 -265 17 -264
rect 39 -262 79 -261
rect 39 -265 79 -264
rect -92 -293 -52 -292
rect 107 -293 108 -253
rect 110 -293 111 -253
rect -92 -296 -52 -295
rect -89 -376 -49 -375
rect -89 -379 -49 -378
rect -20 -376 20 -375
rect -20 -379 20 -378
rect 42 -376 82 -375
rect 42 -379 82 -378
rect -89 -407 -49 -406
rect 110 -407 111 -367
rect 113 -407 114 -367
rect 339 -378 340 -338
rect 342 -378 343 -338
rect 378 -374 379 -334
rect 381 -374 382 -334
rect 411 -368 412 -328
rect 414 -368 415 -328
rect 561 -347 562 -307
rect 564 -347 565 -307
rect 594 -341 595 -301
rect 597 -341 598 -301
rect 670 -336 671 -296
rect 673 -336 674 -296
rect 703 -336 704 -296
rect 706 -336 707 -296
rect 805 -339 806 -299
rect 808 -339 809 -299
rect 838 -333 839 -293
rect 841 -333 842 -293
rect 877 -329 878 -289
rect 880 -329 881 -289
rect -89 -410 -49 -409
<< ndcontact >>
rect 252 670 272 674
rect 252 662 272 666
rect 252 584 272 588
rect 797 624 837 628
rect 851 622 855 642
rect 859 622 863 642
rect 797 616 837 620
rect 252 576 272 580
rect 199 556 203 576
rect 207 556 211 576
rect 308 567 312 587
rect 316 567 320 587
rect 341 567 345 587
rect 349 567 353 587
rect 424 574 464 578
rect 478 572 482 592
rect 486 572 490 592
rect 594 595 634 599
rect 648 593 652 613
rect 656 593 660 613
rect 797 605 837 609
rect 797 597 837 601
rect 594 587 634 591
rect 797 586 837 590
rect 424 566 464 570
rect 594 576 634 580
rect 797 578 837 582
rect 594 568 634 572
rect 797 567 837 571
rect 424 555 464 559
rect 594 557 634 561
rect 797 559 837 563
rect 424 547 464 551
rect 594 549 634 553
rect 797 548 837 552
rect 264 532 284 536
rect 424 536 464 540
rect 594 538 634 542
rect 797 540 837 544
rect 424 528 464 532
rect 594 530 634 534
rect 264 524 284 528
rect 264 446 284 450
rect 264 438 284 442
rect -10 402 10 406
rect 52 402 72 406
rect -10 394 10 398
rect 52 394 72 398
rect 211 418 215 438
rect 219 418 223 438
rect 320 429 324 449
rect 328 429 332 449
rect 353 429 357 449
rect 361 429 365 449
rect 440 432 480 436
rect 494 430 498 450
rect 502 430 506 450
rect 440 424 480 428
rect 610 434 650 438
rect 664 432 668 452
rect 672 432 676 452
rect 610 426 650 430
rect 440 413 480 417
rect 610 415 650 419
rect 1133 433 1153 437
rect 1195 433 1215 437
rect 440 405 480 409
rect 610 407 650 411
rect -106 371 -86 375
rect -36 371 -16 375
rect 26 371 46 375
rect -106 363 -86 367
rect -36 363 -16 367
rect 26 363 46 367
rect 317 394 337 398
rect 317 386 337 390
rect 440 394 480 398
rect 610 396 650 400
rect 440 386 480 390
rect 610 388 650 392
rect 610 378 650 382
rect 686 378 690 398
rect 694 378 698 398
rect 707 378 711 398
rect 715 378 719 398
rect 736 378 740 398
rect 744 378 748 398
rect 769 378 773 398
rect 777 378 781 398
rect 796 378 800 398
rect 804 378 808 398
rect 1133 425 1153 429
rect 1195 425 1215 429
rect 1037 402 1057 406
rect 1107 402 1127 406
rect 1169 402 1189 406
rect 1037 394 1057 398
rect 1107 394 1127 398
rect 1169 394 1189 398
rect 97 345 101 365
rect 105 345 109 365
rect 610 370 650 374
rect 1240 376 1244 396
rect 1248 376 1252 396
rect -11 288 9 292
rect 51 288 71 292
rect -11 280 9 284
rect 51 280 71 284
rect 317 308 337 312
rect 818 350 822 370
rect 826 350 830 370
rect 838 350 842 370
rect 846 350 850 370
rect 859 350 863 370
rect 867 350 871 370
rect 888 350 892 370
rect 896 350 900 370
rect 921 350 925 370
rect 929 350 933 370
rect 948 350 952 370
rect 956 350 960 370
rect 317 300 337 304
rect -107 257 -87 261
rect -37 257 -17 261
rect 25 257 45 261
rect -107 249 -87 253
rect -37 249 -17 253
rect 25 249 45 253
rect 264 280 268 300
rect 272 280 276 300
rect 373 291 377 311
rect 381 291 385 311
rect 406 291 410 311
rect 414 291 418 311
rect 496 271 536 275
rect 550 269 554 289
rect 558 269 562 289
rect 496 263 536 267
rect 317 256 337 260
rect 96 231 100 251
rect 104 231 108 251
rect 317 248 337 252
rect 496 252 536 256
rect 496 244 536 248
rect 593 239 597 259
rect 601 239 605 259
rect 622 239 626 259
rect 630 239 634 259
rect 655 239 659 259
rect 663 239 667 259
rect 682 239 686 259
rect 690 239 694 259
rect 784 261 804 265
rect -8 174 12 178
rect 54 174 74 178
rect -8 166 12 170
rect 54 166 74 170
rect 496 233 536 237
rect 731 234 735 254
rect 739 234 743 254
rect 784 253 804 257
rect 816 233 820 253
rect 824 233 828 253
rect 840 245 844 265
rect 848 245 852 265
rect 873 245 877 265
rect 881 245 885 265
rect 496 225 536 229
rect -104 143 -84 147
rect -34 143 -14 147
rect 28 143 48 147
rect -104 135 -84 139
rect -34 135 -14 139
rect 28 135 48 139
rect 317 170 337 174
rect 317 162 337 166
rect 264 142 268 162
rect 272 142 276 162
rect 373 153 377 173
rect 381 153 385 173
rect 406 153 410 173
rect 414 153 418 173
rect 99 117 103 137
rect 107 117 111 137
rect 610 139 630 143
rect 610 131 630 135
rect -5 60 15 64
rect 57 60 77 64
rect -5 52 15 56
rect 57 52 77 56
rect 264 85 268 105
rect 272 85 276 105
rect 297 85 301 105
rect 305 85 309 105
rect 321 97 325 117
rect 329 97 333 117
rect 345 93 365 97
rect 406 96 410 116
rect 414 96 418 116
rect 450 101 454 121
rect 458 101 462 121
rect 483 101 487 121
rect 491 101 495 121
rect 510 101 514 121
rect 518 101 522 121
rect 345 85 365 89
rect -101 29 -81 33
rect -31 29 -11 33
rect 31 29 51 33
rect -101 21 -81 25
rect -31 21 -11 25
rect 31 21 51 25
rect 1114 113 1134 117
rect 1176 113 1196 117
rect 1114 105 1134 109
rect 1176 105 1196 109
rect 1018 82 1038 86
rect 1088 82 1108 86
rect 1150 82 1170 86
rect 610 53 630 57
rect 1018 74 1038 78
rect 1088 74 1108 78
rect 1150 74 1170 78
rect 1221 56 1225 76
rect 1229 56 1233 76
rect 610 45 630 49
rect 557 25 561 45
rect 565 25 569 45
rect 666 36 670 56
rect 674 36 678 56
rect 699 36 703 56
rect 707 36 711 56
rect 102 3 106 23
rect 110 3 114 23
rect 607 1 627 5
rect 1113 -1 1133 3
rect 1175 -1 1195 3
rect 607 -7 627 -3
rect 1113 -9 1133 -5
rect 1175 -9 1195 -5
rect -6 -58 14 -54
rect 56 -58 76 -54
rect -6 -66 14 -62
rect 56 -66 76 -62
rect 264 -49 268 -29
rect 272 -49 276 -29
rect 297 -49 301 -29
rect 305 -49 309 -29
rect 321 -37 325 -17
rect 329 -37 333 -17
rect 345 -41 365 -37
rect 406 -38 410 -18
rect 414 -38 418 -18
rect 345 -49 365 -45
rect -102 -89 -82 -85
rect -32 -89 -12 -85
rect 30 -89 50 -85
rect -102 -97 -82 -93
rect -32 -97 -12 -93
rect 30 -97 50 -93
rect 101 -115 105 -95
rect 109 -115 113 -95
rect 607 -85 627 -81
rect 1017 -32 1037 -28
rect 1087 -32 1107 -28
rect 1149 -32 1169 -28
rect 1017 -40 1037 -36
rect 1087 -40 1107 -36
rect 1149 -40 1169 -36
rect 1220 -58 1224 -38
rect 1228 -58 1232 -38
rect 607 -93 627 -89
rect 554 -113 558 -93
rect 562 -113 566 -93
rect 663 -102 667 -82
rect 671 -102 675 -82
rect 696 -102 700 -82
rect 704 -102 708 -82
rect 844 -86 864 -82
rect 791 -113 795 -93
rect 799 -113 803 -93
rect 844 -94 864 -90
rect 876 -114 880 -94
rect 884 -114 888 -94
rect 1116 -115 1136 -111
rect 1178 -115 1198 -111
rect 1116 -123 1136 -119
rect 1178 -123 1198 -119
rect 610 -137 630 -133
rect -7 -172 13 -168
rect 55 -172 75 -168
rect -7 -180 13 -176
rect 55 -180 75 -176
rect 610 -145 630 -141
rect 1020 -146 1040 -142
rect 1090 -146 1110 -142
rect 322 -171 326 -151
rect 330 -171 334 -151
rect 1152 -146 1172 -142
rect 346 -175 366 -171
rect 407 -172 411 -152
rect 415 -172 419 -152
rect 1020 -154 1040 -150
rect 1090 -154 1110 -150
rect 1152 -154 1172 -150
rect -103 -203 -83 -199
rect -33 -203 -13 -199
rect 29 -203 49 -199
rect -103 -211 -83 -207
rect -33 -211 -13 -207
rect 29 -211 49 -207
rect 346 -183 366 -179
rect 100 -229 104 -209
rect 108 -229 112 -209
rect 1223 -172 1227 -152
rect 1231 -172 1235 -152
rect 610 -223 630 -219
rect 841 -220 861 -216
rect 610 -231 630 -227
rect 557 -251 561 -231
rect 565 -251 569 -231
rect 788 -247 792 -227
rect 796 -247 800 -227
rect 841 -228 861 -224
rect 873 -248 877 -228
rect 881 -248 885 -228
rect 1119 -229 1139 -225
rect 1181 -229 1201 -225
rect 1119 -237 1139 -233
rect 1181 -237 1201 -233
rect -4 -286 16 -282
rect 58 -286 78 -282
rect -4 -294 16 -290
rect 58 -294 78 -290
rect 1023 -260 1043 -256
rect 1093 -260 1113 -256
rect 1155 -260 1175 -256
rect 1023 -268 1043 -264
rect 1093 -268 1113 -264
rect 1155 -268 1175 -264
rect 610 -275 630 -271
rect 610 -283 630 -279
rect -100 -317 -80 -313
rect -30 -317 -10 -313
rect 32 -317 52 -313
rect -100 -325 -80 -321
rect -30 -325 -10 -321
rect 32 -325 52 -321
rect 322 -305 326 -285
rect 330 -305 334 -285
rect 1226 -286 1230 -266
rect 1234 -286 1238 -266
rect 346 -309 366 -305
rect 407 -306 411 -286
rect 415 -306 419 -286
rect 346 -317 366 -313
rect 103 -343 107 -323
rect 111 -343 115 -323
rect -1 -400 19 -396
rect 61 -400 81 -396
rect -1 -408 19 -404
rect 61 -408 81 -404
rect 610 -361 630 -357
rect 610 -369 630 -365
rect 557 -389 561 -369
rect 565 -389 569 -369
rect 666 -378 670 -358
rect 674 -378 678 -358
rect 699 -378 703 -358
rect 707 -378 711 -358
rect 854 -354 874 -350
rect 801 -381 805 -361
rect 809 -381 813 -361
rect 854 -362 874 -358
rect 886 -382 890 -362
rect 894 -382 898 -362
rect -97 -431 -77 -427
rect -27 -431 -7 -427
rect 35 -431 55 -427
rect -97 -439 -77 -435
rect -27 -439 -7 -435
rect 35 -439 55 -435
rect 106 -457 110 -437
rect 114 -457 118 -437
<< pdcontact >>
rect 199 598 203 638
rect 207 598 211 638
rect 232 604 236 644
rect 240 604 244 644
rect 308 609 312 649
rect 316 609 320 649
rect 341 609 345 649
rect 349 609 353 649
rect 374 614 378 654
rect 382 614 386 654
rect 407 614 411 654
rect 415 614 419 654
rect 440 614 444 654
rect 448 614 452 654
rect 478 614 482 654
rect 486 614 490 654
rect 511 635 515 675
rect 519 635 523 675
rect 544 635 548 675
rect 552 635 556 675
rect 577 635 581 675
rect 585 635 589 675
rect 610 635 614 675
rect 618 635 622 675
rect 648 635 652 675
rect 656 635 660 675
rect 681 664 685 704
rect 689 664 693 704
rect 714 664 718 704
rect 722 664 726 704
rect 747 664 751 704
rect 755 664 759 704
rect 780 664 784 704
rect 788 664 792 704
rect 813 664 817 704
rect 821 664 825 704
rect 851 664 855 704
rect 859 664 863 704
rect 885 532 925 536
rect 732 527 772 531
rect 885 524 925 528
rect 732 519 772 523
rect 211 460 215 500
rect 219 460 223 500
rect 244 466 248 506
rect 252 466 256 506
rect 320 471 324 511
rect 328 471 332 511
rect 353 471 357 511
rect 361 471 365 511
rect 390 472 394 512
rect 398 472 402 512
rect 423 472 427 512
rect 431 472 435 512
rect 456 472 460 512
rect 464 472 468 512
rect 494 472 498 512
rect 502 472 506 512
rect 527 474 531 514
rect 535 474 539 514
rect 560 474 564 514
rect 568 474 572 514
rect 593 474 597 514
rect 601 474 605 514
rect 626 474 630 514
rect 634 474 638 514
rect 664 474 668 514
rect 672 474 676 514
rect 884 499 924 503
rect 731 493 771 497
rect 884 491 924 495
rect 731 485 771 489
rect 883 465 923 469
rect 731 458 771 462
rect -98 427 -58 431
rect -29 427 11 431
rect 33 427 73 431
rect -98 419 -58 423
rect -29 419 11 423
rect 33 419 73 423
rect -98 396 -58 400
rect 97 395 101 435
rect 105 395 109 435
rect 731 450 771 454
rect 731 425 771 429
rect 731 417 771 421
rect 796 420 800 460
rect 804 420 808 460
rect 883 457 923 461
rect 1045 458 1085 462
rect 1114 458 1154 462
rect 1176 458 1216 462
rect 1045 450 1085 454
rect 1114 450 1154 454
rect 1176 450 1216 454
rect 883 430 923 434
rect 883 422 923 426
rect -98 388 -58 392
rect 883 397 923 401
rect 883 389 923 393
rect 948 392 952 432
rect 956 392 960 432
rect 1045 427 1085 431
rect 1240 426 1244 466
rect 1248 426 1252 466
rect 1045 419 1085 423
rect 264 322 268 362
rect 272 322 276 362
rect 297 328 301 368
rect 305 328 309 368
rect 373 333 377 373
rect 381 333 385 373
rect 406 333 410 373
rect 414 333 418 373
rect 617 354 657 358
rect -99 313 -59 317
rect -30 313 10 317
rect 32 313 72 317
rect -99 305 -59 309
rect -30 305 10 309
rect 32 305 72 309
rect -99 282 -59 286
rect 96 281 100 321
rect 104 281 108 321
rect 446 311 450 351
rect 454 311 458 351
rect 479 311 483 351
rect 487 311 491 351
rect 512 311 516 351
rect 520 311 524 351
rect 550 311 554 351
rect 558 311 562 351
rect 617 346 657 350
rect 617 319 657 323
rect 617 311 657 315
rect -99 274 -59 278
rect 617 286 657 290
rect 617 278 657 282
rect 682 281 686 321
rect 690 281 694 321
rect 731 276 735 316
rect 739 276 743 316
rect 764 282 768 322
rect 772 282 776 322
rect 803 286 807 326
rect 811 286 815 326
rect 840 287 844 327
rect 848 287 852 327
rect 873 287 877 327
rect 881 287 885 327
rect -96 199 -56 203
rect -27 199 13 203
rect 35 199 75 203
rect -96 191 -56 195
rect -27 191 13 195
rect 35 191 75 195
rect -96 168 -56 172
rect 99 167 103 207
rect 107 167 111 207
rect 264 184 268 224
rect 272 184 276 224
rect 297 190 301 230
rect 305 190 309 230
rect 373 195 377 235
rect 381 195 385 235
rect 406 195 410 235
rect 414 195 418 235
rect -96 160 -56 164
rect 445 181 485 185
rect 445 173 485 177
rect 445 148 485 152
rect 445 140 485 144
rect 510 143 514 183
rect 518 143 522 183
rect 1026 138 1066 142
rect 1095 138 1135 142
rect 1157 138 1197 142
rect 1026 130 1066 134
rect 1095 130 1135 134
rect 1157 130 1197 134
rect -93 85 -53 89
rect -24 85 16 89
rect 38 85 78 89
rect -93 77 -53 81
rect -24 77 16 81
rect 38 77 78 81
rect -93 54 -53 58
rect 102 53 106 93
rect 110 53 114 93
rect -93 46 -53 50
rect 264 23 268 63
rect 272 23 276 63
rect 297 23 301 63
rect 305 23 309 63
rect 334 24 338 64
rect 342 24 346 64
rect 373 28 377 68
rect 381 28 385 68
rect 406 34 410 74
rect 414 34 418 74
rect 557 67 561 107
rect 565 67 569 107
rect 590 73 594 113
rect 598 73 602 113
rect 666 78 670 118
rect 674 78 678 118
rect 699 78 703 118
rect 707 78 711 118
rect 1026 107 1066 111
rect 1221 106 1225 146
rect 1229 106 1233 146
rect 1026 99 1066 103
rect 1025 24 1065 28
rect 1094 24 1134 28
rect 1156 24 1196 28
rect 1025 16 1065 20
rect 1094 16 1134 20
rect 1156 16 1196 20
rect 1025 -7 1065 -3
rect 1220 -8 1224 32
rect 1228 -8 1232 32
rect 1025 -15 1065 -11
rect -94 -33 -54 -29
rect -25 -33 15 -29
rect 37 -33 77 -29
rect -94 -41 -54 -37
rect -25 -41 15 -37
rect 37 -41 77 -37
rect -94 -64 -54 -60
rect 101 -65 105 -25
rect 109 -65 113 -25
rect -94 -72 -54 -68
rect 264 -111 268 -71
rect 272 -111 276 -71
rect 297 -111 301 -71
rect 305 -111 309 -71
rect 334 -110 338 -70
rect 342 -110 346 -70
rect 373 -106 377 -66
rect 381 -106 385 -66
rect 406 -100 410 -60
rect 414 -100 418 -60
rect 554 -71 558 -31
rect 562 -71 566 -31
rect 587 -65 591 -25
rect 595 -65 599 -25
rect 663 -60 667 -20
rect 671 -60 675 -20
rect 696 -60 700 -20
rect 704 -60 708 -20
rect 791 -71 795 -31
rect 799 -71 803 -31
rect 824 -65 828 -25
rect 832 -65 836 -25
rect 863 -61 867 -21
rect 871 -61 875 -21
rect 1028 -90 1068 -86
rect 1097 -90 1137 -86
rect 1159 -90 1199 -86
rect 1028 -98 1068 -94
rect 1097 -98 1137 -94
rect 1159 -98 1199 -94
rect 1028 -121 1068 -117
rect 1223 -122 1227 -82
rect 1231 -122 1235 -82
rect 1028 -129 1068 -125
rect -95 -147 -55 -143
rect -26 -147 14 -143
rect 36 -147 76 -143
rect -95 -155 -55 -151
rect -26 -155 14 -151
rect 36 -155 76 -151
rect -95 -178 -55 -174
rect 100 -179 104 -139
rect 108 -179 112 -139
rect -95 -186 -55 -182
rect 335 -244 339 -204
rect 343 -244 347 -204
rect 374 -240 378 -200
rect 382 -240 386 -200
rect 407 -234 411 -194
rect 415 -234 419 -194
rect 557 -209 561 -169
rect 565 -209 569 -169
rect 590 -203 594 -163
rect 598 -203 602 -163
rect 788 -205 792 -165
rect 796 -205 800 -165
rect 821 -199 825 -159
rect 829 -199 833 -159
rect 860 -195 864 -155
rect 868 -195 872 -155
rect 1031 -204 1071 -200
rect 1100 -204 1140 -200
rect 1162 -204 1202 -200
rect 1031 -212 1071 -208
rect 1100 -212 1140 -208
rect 1162 -212 1202 -208
rect 1031 -235 1071 -231
rect 1226 -236 1230 -196
rect 1234 -236 1238 -196
rect 1031 -243 1071 -239
rect -92 -261 -52 -257
rect -23 -261 17 -257
rect 39 -261 79 -257
rect -92 -269 -52 -265
rect -23 -269 17 -265
rect 39 -269 79 -265
rect -92 -292 -52 -288
rect 103 -293 107 -253
rect 111 -293 115 -253
rect -92 -300 -52 -296
rect -89 -375 -49 -371
rect -20 -375 20 -371
rect 42 -375 82 -371
rect -89 -383 -49 -379
rect -20 -383 20 -379
rect 42 -383 82 -379
rect -89 -406 -49 -402
rect 106 -407 110 -367
rect 114 -407 118 -367
rect 335 -378 339 -338
rect 343 -378 347 -338
rect 374 -374 378 -334
rect 382 -374 386 -334
rect 407 -368 411 -328
rect 415 -368 419 -328
rect 557 -347 561 -307
rect 565 -347 569 -307
rect 590 -341 594 -301
rect 598 -341 602 -301
rect 666 -336 670 -296
rect 674 -336 678 -296
rect 699 -336 703 -296
rect 707 -336 711 -296
rect 801 -339 805 -299
rect 809 -339 813 -299
rect 834 -333 838 -293
rect 842 -333 846 -293
rect 873 -329 877 -289
rect 881 -329 885 -289
rect -89 -414 -49 -410
<< polysilicon >>
rect 686 704 688 707
rect 719 704 721 707
rect 752 704 754 707
rect 785 704 787 707
rect 818 704 820 707
rect 856 704 858 707
rect 516 675 518 678
rect 549 675 551 678
rect 582 675 584 678
rect 615 675 617 678
rect 653 675 655 678
rect 249 667 252 669
rect 272 667 275 669
rect 379 654 381 657
rect 412 654 414 657
rect 445 654 447 657
rect 483 654 485 657
rect 313 649 315 652
rect 346 649 348 652
rect 237 644 239 647
rect 204 638 206 641
rect 686 651 688 664
rect 719 651 721 664
rect 752 651 754 664
rect 785 651 787 664
rect 818 651 820 664
rect 856 642 858 664
rect 516 622 518 635
rect 549 622 551 635
rect 582 622 584 635
rect 615 622 617 635
rect 204 576 206 598
rect 237 592 239 604
rect 313 587 315 609
rect 346 587 348 609
rect 379 601 381 614
rect 412 601 414 614
rect 445 601 447 614
rect 483 592 485 614
rect 653 613 655 635
rect 794 621 797 623
rect 837 621 840 623
rect 856 619 858 622
rect 244 581 252 583
rect 272 581 275 583
rect 421 571 424 573
rect 464 571 467 573
rect 591 592 594 594
rect 634 592 637 594
rect 794 602 797 604
rect 837 602 840 604
rect 653 590 655 593
rect 794 583 797 585
rect 837 583 840 585
rect 313 564 315 567
rect 346 564 348 567
rect 483 569 485 572
rect 591 573 594 575
rect 634 573 637 575
rect 794 564 797 566
rect 837 564 840 566
rect 204 553 206 556
rect 421 552 424 554
rect 464 552 467 554
rect 591 554 594 556
rect 634 554 637 556
rect 794 545 797 547
rect 837 545 840 547
rect 421 533 424 535
rect 464 533 467 535
rect 591 535 594 537
rect 634 535 637 537
rect 261 529 264 531
rect 284 529 287 531
rect 882 529 885 531
rect 925 529 936 531
rect 729 524 732 526
rect 772 524 783 526
rect 325 511 327 514
rect 358 511 360 514
rect 395 512 397 515
rect 428 512 430 515
rect 461 512 463 515
rect 499 512 501 515
rect 532 514 534 517
rect 565 514 567 517
rect 598 514 600 517
rect 631 514 633 517
rect 669 514 671 517
rect 249 506 251 509
rect 216 500 218 503
rect 881 496 884 498
rect 924 496 935 498
rect 728 490 731 492
rect 771 490 782 492
rect 216 438 218 460
rect 249 454 251 466
rect 325 449 327 471
rect 358 449 360 471
rect 395 459 397 472
rect 428 459 430 472
rect 461 459 463 472
rect 499 450 501 472
rect 532 461 534 474
rect 565 461 567 474
rect 598 461 600 474
rect 631 461 633 474
rect 669 452 671 474
rect 1245 466 1247 469
rect 801 460 803 463
rect 880 462 883 464
rect 923 462 934 464
rect 728 455 731 457
rect 771 455 782 457
rect 256 443 264 445
rect 284 443 287 445
rect 102 435 104 438
rect -108 424 -98 426
rect -58 424 -55 426
rect -39 424 -29 426
rect 11 424 14 426
rect 24 424 33 426
rect 73 424 76 426
rect -13 399 -10 401
rect 10 399 13 401
rect 49 399 52 401
rect 72 399 75 401
rect -108 393 -98 395
rect -58 393 -55 395
rect 325 426 327 429
rect 358 426 360 429
rect 437 429 440 431
rect 480 429 483 431
rect 499 427 501 430
rect 607 431 610 433
rect 650 431 653 433
rect 669 429 671 432
rect 728 422 731 424
rect 771 422 777 424
rect 216 415 218 418
rect 437 410 440 412
rect 480 410 483 412
rect 775 418 777 422
rect 1035 455 1045 457
rect 1085 455 1088 457
rect 1104 455 1114 457
rect 1154 455 1157 457
rect 1167 455 1176 457
rect 1216 455 1219 457
rect 953 432 955 435
rect 880 427 883 429
rect 923 427 934 429
rect 607 412 610 414
rect 650 412 653 414
rect -109 368 -106 370
rect -86 368 -83 370
rect -39 368 -36 370
rect -16 368 -13 370
rect 23 368 26 370
rect 46 368 49 370
rect 102 365 104 395
rect 314 391 317 393
rect 337 391 340 393
rect 437 391 440 393
rect 480 391 483 393
rect 691 398 693 401
rect 712 398 714 401
rect 741 398 743 401
rect 774 398 776 401
rect 801 398 803 420
rect 607 393 610 395
rect 650 393 653 395
rect 378 373 380 376
rect 411 373 413 376
rect 880 394 883 396
rect 923 394 929 396
rect 927 390 929 394
rect 1130 430 1133 432
rect 1153 430 1156 432
rect 1192 430 1195 432
rect 1215 430 1218 432
rect 1035 424 1045 426
rect 1085 424 1088 426
rect 1034 399 1037 401
rect 1057 399 1060 401
rect 1104 399 1107 401
rect 1127 399 1130 401
rect 1166 399 1169 401
rect 1189 399 1192 401
rect 1245 396 1247 426
rect 607 375 610 377
rect 650 375 653 377
rect 691 375 693 378
rect 712 375 714 378
rect 741 375 743 378
rect 774 375 776 378
rect 801 375 803 378
rect 302 368 304 371
rect 269 362 271 365
rect 102 342 104 345
rect 101 321 103 324
rect 823 370 825 373
rect 843 370 845 373
rect 864 370 866 373
rect 893 370 895 373
rect 926 370 928 373
rect 953 370 955 392
rect 1245 373 1247 376
rect 451 351 453 354
rect 484 351 486 354
rect 517 351 519 354
rect 555 351 557 354
rect -109 310 -99 312
rect -59 310 -56 312
rect -40 310 -30 312
rect 10 310 13 312
rect 23 310 32 312
rect 72 310 75 312
rect -14 285 -11 287
rect 9 285 12 287
rect 48 285 51 287
rect 71 285 74 287
rect -109 279 -99 281
rect -59 279 -56 281
rect 269 300 271 322
rect 302 316 304 328
rect 378 311 380 333
rect 411 311 413 333
rect 614 351 617 353
rect 657 351 668 353
rect 823 347 825 350
rect 843 347 845 350
rect 864 347 866 350
rect 893 347 895 350
rect 926 347 928 350
rect 953 347 955 350
rect 808 326 810 329
rect 845 327 847 330
rect 878 327 880 330
rect 687 321 689 324
rect 769 322 771 325
rect 614 316 617 318
rect 657 316 668 318
rect 309 305 317 307
rect 337 305 340 307
rect -110 254 -107 256
rect -87 254 -84 256
rect -40 254 -37 256
rect -17 254 -14 256
rect 22 254 25 256
rect 45 254 48 256
rect 101 251 103 281
rect 451 298 453 311
rect 484 298 486 311
rect 517 298 519 311
rect 378 288 380 291
rect 411 288 413 291
rect 555 289 557 311
rect 269 277 271 280
rect 493 268 496 270
rect 536 268 539 270
rect 614 283 617 285
rect 657 283 663 285
rect 661 279 663 283
rect 736 316 738 319
rect 555 266 557 269
rect 598 259 600 262
rect 627 259 629 262
rect 660 259 662 262
rect 687 259 689 281
rect 808 283 810 286
rect 769 276 771 282
rect 314 253 317 255
rect 337 253 340 255
rect 493 249 496 251
rect 536 249 539 251
rect 736 254 738 276
rect 845 265 847 287
rect 878 265 880 287
rect 776 258 784 260
rect 804 258 807 260
rect 378 235 380 238
rect 411 235 413 238
rect 101 228 103 231
rect 302 230 304 233
rect 269 224 271 227
rect 104 207 106 210
rect -106 196 -96 198
rect -56 196 -53 198
rect -37 196 -27 198
rect 13 196 16 198
rect 26 196 35 198
rect 75 196 78 198
rect -11 171 -8 173
rect 12 171 15 173
rect 51 171 54 173
rect 74 171 77 173
rect -106 165 -96 167
rect -56 165 -53 167
rect 598 236 600 239
rect 627 236 629 239
rect 660 236 662 239
rect 687 236 689 239
rect 821 253 823 257
rect 493 230 496 232
rect 536 230 539 232
rect 736 231 738 234
rect 845 242 847 245
rect 878 242 880 245
rect 821 230 823 233
rect -107 140 -104 142
rect -84 140 -81 142
rect -37 140 -34 142
rect -14 140 -11 142
rect 25 140 28 142
rect 48 140 51 142
rect 104 137 106 167
rect 269 162 271 184
rect 302 178 304 190
rect 378 173 380 195
rect 411 173 413 195
rect 515 183 517 186
rect 442 178 445 180
rect 485 178 496 180
rect 309 167 317 169
rect 337 167 340 169
rect 378 150 380 153
rect 411 150 413 153
rect 442 145 445 147
rect 485 145 491 147
rect 269 139 271 142
rect 489 141 491 145
rect 1226 146 1228 149
rect 455 121 457 124
rect 488 121 490 124
rect 515 121 517 143
rect 607 136 610 138
rect 630 136 633 138
rect 1016 135 1026 137
rect 1066 135 1069 137
rect 1085 135 1095 137
rect 1135 135 1138 137
rect 1148 135 1157 137
rect 1197 135 1200 137
rect 326 117 328 120
rect 104 114 106 117
rect 269 105 271 108
rect 302 105 304 108
rect 107 93 109 96
rect -103 82 -93 84
rect -53 82 -50 84
rect -34 82 -24 84
rect 16 82 19 84
rect 29 82 38 84
rect 78 82 81 84
rect -8 57 -5 59
rect 15 57 18 59
rect 54 57 57 59
rect 77 57 80 59
rect -103 51 -93 53
rect -53 51 -50 53
rect 411 116 413 119
rect 326 93 328 97
rect 671 118 673 121
rect 704 118 706 121
rect 595 113 597 116
rect 562 107 564 110
rect 455 98 457 101
rect 488 98 490 101
rect 515 98 517 101
rect 342 90 345 92
rect 365 90 373 92
rect 269 63 271 85
rect 302 63 304 85
rect 411 74 413 96
rect 378 68 380 74
rect 339 64 341 67
rect -104 26 -101 28
rect -81 26 -78 28
rect -34 26 -31 28
rect -11 26 -8 28
rect 28 26 31 28
rect 51 26 54 28
rect 107 23 109 53
rect 1111 110 1114 112
rect 1134 110 1137 112
rect 1173 110 1176 112
rect 1196 110 1199 112
rect 1016 104 1026 106
rect 1066 104 1069 106
rect 1015 79 1018 81
rect 1038 79 1041 81
rect 1085 79 1088 81
rect 1108 79 1111 81
rect 1147 79 1150 81
rect 1170 79 1173 81
rect 562 45 564 67
rect 595 61 597 73
rect 671 56 673 78
rect 704 56 706 78
rect 1226 76 1228 106
rect 602 50 610 52
rect 630 50 633 52
rect 411 31 413 34
rect 378 25 380 28
rect 1226 53 1228 56
rect 671 33 673 36
rect 704 33 706 36
rect 1225 32 1227 35
rect 269 20 271 23
rect 302 20 304 23
rect 339 21 341 24
rect 562 22 564 25
rect 1015 21 1025 23
rect 1065 21 1068 23
rect 1084 21 1094 23
rect 1134 21 1137 23
rect 1147 21 1156 23
rect 1196 21 1199 23
rect 107 0 109 3
rect 604 -2 607 0
rect 627 -2 630 0
rect 1110 -4 1113 -2
rect 1133 -4 1136 -2
rect 1172 -4 1175 -2
rect 1195 -4 1198 -2
rect 1015 -10 1025 -8
rect 1065 -10 1068 -8
rect 326 -17 328 -14
rect 106 -25 108 -22
rect -104 -36 -94 -34
rect -54 -36 -51 -34
rect -35 -36 -25 -34
rect 15 -36 18 -34
rect 28 -36 37 -34
rect 77 -36 80 -34
rect -9 -61 -6 -59
rect 14 -61 17 -59
rect 53 -61 56 -59
rect 76 -61 79 -59
rect -104 -67 -94 -65
rect -54 -67 -51 -65
rect 269 -29 271 -26
rect 302 -29 304 -26
rect 411 -18 413 -15
rect 326 -41 328 -37
rect 668 -20 670 -17
rect 701 -20 703 -17
rect 592 -25 594 -22
rect 559 -31 561 -28
rect 342 -44 345 -42
rect 365 -44 373 -42
rect -105 -92 -102 -90
rect -82 -92 -79 -90
rect -35 -92 -32 -90
rect -12 -92 -9 -90
rect 27 -92 30 -90
rect 50 -92 53 -90
rect 106 -95 108 -65
rect 269 -71 271 -49
rect 302 -71 304 -49
rect 411 -60 413 -38
rect 378 -66 380 -60
rect 339 -70 341 -67
rect 868 -21 870 -18
rect 829 -25 831 -22
rect 796 -31 798 -28
rect 559 -93 561 -71
rect 592 -77 594 -65
rect 668 -82 670 -60
rect 701 -82 703 -60
rect 1014 -35 1017 -33
rect 1037 -35 1040 -33
rect 1084 -35 1087 -33
rect 1107 -35 1110 -33
rect 1146 -35 1149 -33
rect 1169 -35 1172 -33
rect 1225 -38 1227 -8
rect 1225 -61 1227 -58
rect 868 -64 870 -61
rect 829 -71 831 -65
rect 599 -88 607 -86
rect 627 -88 630 -86
rect 411 -103 413 -100
rect 378 -109 380 -106
rect 269 -114 271 -111
rect 302 -114 304 -111
rect 339 -113 341 -110
rect 796 -93 798 -71
rect 1228 -82 1230 -79
rect 836 -89 844 -87
rect 864 -89 867 -87
rect 668 -105 670 -102
rect 701 -105 703 -102
rect 881 -94 883 -90
rect 1018 -93 1028 -91
rect 1068 -93 1071 -91
rect 1087 -93 1097 -91
rect 1137 -93 1140 -91
rect 1150 -93 1159 -91
rect 1199 -93 1202 -91
rect 106 -118 108 -115
rect 559 -116 561 -113
rect 796 -116 798 -113
rect 881 -117 883 -114
rect 1113 -118 1116 -116
rect 1136 -118 1139 -116
rect 1175 -118 1178 -116
rect 1198 -118 1201 -116
rect 1018 -124 1028 -122
rect 1068 -124 1071 -122
rect 105 -139 107 -136
rect -105 -150 -95 -148
rect -55 -150 -52 -148
rect -36 -150 -26 -148
rect 14 -150 17 -148
rect 27 -150 36 -148
rect 76 -150 79 -148
rect -10 -175 -7 -173
rect 13 -175 16 -173
rect 52 -175 55 -173
rect 75 -175 78 -173
rect -105 -181 -95 -179
rect -55 -181 -52 -179
rect 607 -140 610 -138
rect 630 -140 633 -138
rect 327 -151 329 -148
rect 412 -152 414 -149
rect 1017 -149 1020 -147
rect 1040 -149 1043 -147
rect 1087 -149 1090 -147
rect 1110 -149 1113 -147
rect 1149 -149 1152 -147
rect 1172 -149 1175 -147
rect 327 -175 329 -171
rect 865 -155 867 -152
rect 1228 -152 1230 -122
rect 826 -159 828 -156
rect 595 -163 597 -160
rect 562 -169 564 -166
rect -106 -206 -103 -204
rect -83 -206 -80 -204
rect -36 -206 -33 -204
rect -13 -206 -10 -204
rect 26 -206 29 -204
rect 49 -206 52 -204
rect 105 -209 107 -179
rect 343 -178 346 -176
rect 366 -178 374 -176
rect 412 -194 414 -172
rect 379 -200 381 -194
rect 340 -204 342 -201
rect 105 -232 107 -229
rect 793 -165 795 -162
rect 562 -231 564 -209
rect 595 -215 597 -203
rect 1228 -175 1230 -172
rect 865 -198 867 -195
rect 1231 -196 1233 -193
rect 826 -205 828 -199
rect 602 -226 610 -224
rect 630 -226 633 -224
rect 793 -227 795 -205
rect 1021 -207 1031 -205
rect 1071 -207 1074 -205
rect 1090 -207 1100 -205
rect 1140 -207 1143 -205
rect 1153 -207 1162 -205
rect 1202 -207 1205 -205
rect 833 -223 841 -221
rect 861 -223 864 -221
rect 412 -237 414 -234
rect 379 -243 381 -240
rect 340 -247 342 -244
rect 108 -253 110 -250
rect 878 -228 880 -224
rect 793 -250 795 -247
rect 1116 -232 1119 -230
rect 1139 -232 1142 -230
rect 1178 -232 1181 -230
rect 1201 -232 1204 -230
rect 1021 -238 1031 -236
rect 1071 -238 1074 -236
rect 878 -251 880 -248
rect -102 -264 -92 -262
rect -52 -264 -49 -262
rect -33 -264 -23 -262
rect 17 -264 20 -262
rect 30 -264 39 -262
rect 79 -264 82 -262
rect -7 -289 -4 -287
rect 16 -289 19 -287
rect 55 -289 58 -287
rect 78 -289 81 -287
rect -102 -295 -92 -293
rect -52 -295 -49 -293
rect 562 -254 564 -251
rect 1020 -263 1023 -261
rect 1043 -263 1046 -261
rect 1090 -263 1093 -261
rect 1113 -263 1116 -261
rect 1152 -263 1155 -261
rect 1175 -263 1178 -261
rect 1231 -266 1233 -236
rect 607 -278 610 -276
rect 630 -278 633 -276
rect 327 -285 329 -282
rect -103 -320 -100 -318
rect -80 -320 -77 -318
rect -33 -320 -30 -318
rect -10 -320 -7 -318
rect 29 -320 32 -318
rect 52 -320 55 -318
rect 108 -323 110 -293
rect 412 -286 414 -283
rect 327 -309 329 -305
rect 878 -289 880 -286
rect 1231 -289 1233 -286
rect 839 -293 841 -290
rect 671 -296 673 -293
rect 704 -296 706 -293
rect 595 -301 597 -298
rect 343 -312 346 -310
rect 366 -312 374 -310
rect 412 -328 414 -306
rect 562 -307 564 -304
rect 379 -334 381 -328
rect 340 -338 342 -335
rect 108 -346 110 -343
rect 111 -367 113 -364
rect -99 -378 -89 -376
rect -49 -378 -46 -376
rect -30 -378 -20 -376
rect 20 -378 23 -376
rect 33 -378 42 -376
rect 82 -378 85 -376
rect -4 -403 -1 -401
rect 19 -403 22 -401
rect 58 -403 61 -401
rect 81 -403 84 -401
rect -99 -409 -89 -407
rect -49 -409 -46 -407
rect 806 -299 808 -296
rect 412 -371 414 -368
rect 562 -369 564 -347
rect 595 -353 597 -341
rect 671 -358 673 -336
rect 704 -358 706 -336
rect 878 -332 880 -329
rect 839 -339 841 -333
rect 602 -364 610 -362
rect 630 -364 633 -362
rect 379 -377 381 -374
rect 340 -381 342 -378
rect 806 -361 808 -339
rect 846 -357 854 -355
rect 874 -357 877 -355
rect 671 -381 673 -378
rect 704 -381 706 -378
rect 891 -362 893 -358
rect 806 -384 808 -381
rect 891 -385 893 -382
rect 562 -392 564 -389
rect -100 -434 -97 -432
rect -77 -434 -74 -432
rect -30 -434 -27 -432
rect -7 -434 -4 -432
rect 32 -434 35 -432
rect 55 -434 58 -432
rect 111 -437 113 -407
rect 111 -460 113 -457
<< polycontact >>
rect 245 666 249 670
rect 685 647 689 651
rect 718 647 722 651
rect 751 647 755 651
rect 784 647 788 651
rect 817 647 821 651
rect 852 646 856 650
rect 515 618 519 622
rect 548 618 552 622
rect 581 618 585 622
rect 614 618 618 622
rect 649 617 653 621
rect 200 580 204 584
rect 236 588 240 592
rect 309 591 313 595
rect 342 591 346 595
rect 378 597 382 601
rect 411 597 415 601
rect 444 597 448 601
rect 479 596 483 600
rect 788 619 794 625
rect 240 580 244 584
rect 415 569 421 575
rect 585 590 591 596
rect 788 600 794 606
rect 788 581 794 587
rect 585 571 591 577
rect 788 562 794 568
rect 415 550 421 556
rect 585 552 591 558
rect 788 543 794 549
rect 257 528 261 532
rect 415 531 421 537
rect 585 533 591 539
rect 878 528 882 532
rect 725 523 729 527
rect 877 495 881 499
rect 724 489 728 493
rect 212 442 216 446
rect 248 450 252 454
rect 321 453 325 457
rect 354 453 358 457
rect 394 455 398 459
rect 427 455 431 459
rect 460 455 464 459
rect 495 454 499 458
rect 531 457 535 461
rect 564 457 568 461
rect 597 457 601 461
rect 630 457 634 461
rect 665 456 669 460
rect 876 461 880 465
rect 724 454 728 458
rect 252 442 256 446
rect -112 423 -108 427
rect -43 423 -39 427
rect 20 423 24 427
rect -17 398 -13 402
rect 45 398 49 402
rect -112 392 -108 396
rect 431 427 437 433
rect 601 429 607 435
rect 431 408 437 414
rect 601 410 607 416
rect 1031 454 1035 458
rect 1100 454 1104 458
rect 1163 454 1167 458
rect 876 426 880 430
rect 774 414 778 418
rect 690 401 694 405
rect 711 401 715 405
rect 740 401 744 405
rect 774 401 778 405
rect 797 402 801 406
rect -113 367 -109 371
rect -43 367 -39 371
rect 19 368 23 372
rect 98 369 102 373
rect 310 390 314 394
rect 431 389 437 395
rect 601 391 607 397
rect 601 373 607 379
rect 1126 429 1130 433
rect 1188 429 1192 433
rect 1031 423 1035 427
rect 1030 398 1034 402
rect 1100 398 1104 402
rect 1162 399 1166 403
rect 1241 400 1245 404
rect 926 386 930 390
rect 822 373 826 377
rect 842 373 846 377
rect 863 373 867 377
rect 892 373 896 377
rect 926 373 930 377
rect 949 374 953 378
rect -113 309 -109 313
rect -44 309 -40 313
rect 19 309 23 313
rect -18 284 -14 288
rect 44 284 48 288
rect -113 278 -109 282
rect 265 304 269 308
rect 301 312 305 316
rect 374 315 378 319
rect 407 315 411 319
rect 610 350 614 354
rect 768 325 772 329
rect 610 315 614 319
rect 305 304 309 308
rect -114 253 -110 257
rect -44 253 -40 257
rect 18 254 22 258
rect 97 255 101 259
rect 450 294 454 298
rect 483 294 487 298
rect 516 294 520 298
rect 551 293 555 297
rect 487 266 493 272
rect 660 275 664 279
rect 597 262 601 266
rect 626 262 630 266
rect 660 262 664 266
rect 683 263 687 267
rect 806 278 812 283
rect 310 252 314 256
rect 487 247 493 253
rect 732 258 736 262
rect 841 269 845 273
rect 874 269 878 273
rect 772 257 776 261
rect 819 257 825 262
rect -110 195 -106 199
rect -41 195 -37 199
rect 22 195 26 199
rect -15 170 -11 174
rect 47 170 51 174
rect -110 164 -106 168
rect 487 228 493 234
rect -111 139 -107 143
rect -41 139 -37 143
rect 21 140 25 144
rect 100 141 104 145
rect 265 166 269 170
rect 301 174 305 178
rect 374 177 378 181
rect 407 177 411 181
rect 438 177 442 181
rect 305 166 309 170
rect 488 137 492 141
rect 454 124 458 128
rect 488 124 492 128
rect 511 125 515 129
rect 603 135 607 139
rect 1012 134 1016 138
rect 1081 134 1085 138
rect 1144 134 1148 138
rect -107 81 -103 85
rect -38 81 -34 85
rect 25 81 29 85
rect -12 56 -8 60
rect 50 56 54 60
rect -107 50 -103 54
rect 324 88 330 93
rect 373 89 377 93
rect 271 77 275 81
rect 304 77 308 81
rect 413 88 417 92
rect 337 67 343 72
rect -108 25 -104 29
rect -38 25 -34 29
rect 24 26 28 30
rect 103 27 107 31
rect 1107 109 1111 113
rect 1169 109 1173 113
rect 1012 103 1016 107
rect 1011 78 1015 82
rect 1081 78 1085 82
rect 1143 79 1147 83
rect 1222 80 1226 84
rect 558 49 562 53
rect 594 57 598 61
rect 667 60 671 64
rect 700 60 704 64
rect 598 49 602 53
rect 377 21 381 25
rect 1011 20 1015 24
rect 1080 20 1084 24
rect 1143 20 1147 24
rect 600 -3 604 1
rect 1106 -5 1110 -1
rect 1168 -5 1172 -1
rect 1011 -11 1015 -7
rect -108 -37 -104 -33
rect -39 -37 -35 -33
rect 24 -37 28 -33
rect -13 -62 -9 -58
rect 49 -62 53 -58
rect -108 -68 -104 -64
rect 324 -46 330 -41
rect 373 -45 377 -41
rect -109 -93 -105 -89
rect -39 -93 -35 -89
rect 23 -92 27 -88
rect 102 -91 106 -87
rect 271 -57 275 -53
rect 304 -57 308 -53
rect 413 -46 417 -42
rect 337 -67 343 -62
rect 828 -22 832 -18
rect 555 -89 559 -85
rect 591 -81 595 -77
rect 664 -78 668 -74
rect 697 -78 701 -74
rect 1010 -36 1014 -32
rect 1080 -36 1084 -32
rect 1142 -35 1146 -31
rect 1221 -34 1225 -30
rect 866 -69 872 -64
rect 595 -89 599 -85
rect 377 -113 381 -109
rect 792 -89 796 -85
rect 832 -90 836 -86
rect 879 -90 885 -85
rect 1014 -94 1018 -90
rect 1083 -94 1087 -90
rect 1146 -94 1150 -90
rect 1109 -119 1113 -115
rect 1171 -119 1175 -115
rect 1014 -125 1018 -121
rect -109 -151 -105 -147
rect -40 -151 -36 -147
rect 23 -151 27 -147
rect -14 -176 -10 -172
rect 48 -176 52 -172
rect -109 -182 -105 -178
rect 603 -141 607 -137
rect 1013 -150 1017 -146
rect 1083 -150 1087 -146
rect 1145 -149 1149 -145
rect 1224 -148 1228 -144
rect 825 -156 829 -152
rect -110 -207 -106 -203
rect -40 -207 -36 -203
rect 22 -206 26 -202
rect 101 -205 105 -201
rect 325 -180 331 -175
rect 374 -179 378 -175
rect 414 -180 418 -176
rect 338 -201 344 -196
rect 558 -227 562 -223
rect 863 -203 869 -198
rect 594 -219 598 -215
rect 789 -223 793 -219
rect 598 -227 602 -223
rect 1017 -208 1021 -204
rect 1086 -208 1090 -204
rect 1149 -208 1153 -204
rect 829 -224 833 -220
rect 876 -224 882 -219
rect 378 -247 382 -243
rect 1112 -233 1116 -229
rect 1174 -233 1178 -229
rect 1017 -239 1021 -235
rect -106 -265 -102 -261
rect -37 -265 -33 -261
rect 26 -265 30 -261
rect -11 -290 -7 -286
rect 51 -290 55 -286
rect -106 -296 -102 -292
rect 1016 -264 1020 -260
rect 1086 -264 1090 -260
rect 1148 -263 1152 -259
rect 1227 -262 1231 -258
rect 603 -279 607 -275
rect -107 -321 -103 -317
rect -37 -321 -33 -317
rect 25 -320 29 -316
rect 104 -319 108 -315
rect 838 -290 842 -286
rect 325 -314 331 -309
rect 374 -313 378 -309
rect 414 -314 418 -310
rect 338 -335 344 -330
rect -103 -379 -99 -375
rect -34 -379 -30 -375
rect 29 -379 33 -375
rect -8 -404 -4 -400
rect 54 -404 58 -400
rect -103 -410 -99 -406
rect 558 -365 562 -361
rect 594 -357 598 -353
rect 667 -354 671 -350
rect 700 -354 704 -350
rect 876 -337 882 -332
rect 802 -357 806 -353
rect 598 -365 602 -361
rect 378 -381 382 -377
rect 842 -358 846 -354
rect 889 -358 895 -353
rect -104 -435 -100 -431
rect -34 -435 -30 -431
rect 28 -434 32 -430
rect 107 -433 111 -429
<< metal1 >>
rect 663 714 869 717
rect 663 713 699 714
rect 663 688 666 713
rect 675 710 699 713
rect 708 710 732 714
rect 741 710 765 714
rect 774 710 798 714
rect 807 710 831 714
rect 845 710 869 714
rect 493 685 666 688
rect 493 684 529 685
rect 272 670 285 674
rect 185 666 245 670
rect 185 584 190 666
rect 268 653 272 662
rect 193 644 217 651
rect 226 650 272 653
rect 232 644 236 650
rect 199 638 203 644
rect 207 584 211 598
rect 240 599 244 604
rect 279 599 285 670
rect 493 667 496 684
rect 505 681 529 684
rect 538 681 562 685
rect 571 681 595 685
rect 604 681 628 685
rect 642 681 666 685
rect 681 704 685 710
rect 714 704 718 710
rect 747 704 751 710
rect 780 704 784 710
rect 813 704 817 710
rect 851 704 855 710
rect 356 664 496 667
rect 356 663 392 664
rect 356 662 359 663
rect 302 655 359 662
rect 368 660 392 663
rect 401 660 425 664
rect 434 660 458 664
rect 472 660 496 664
rect 511 675 515 681
rect 544 675 548 681
rect 577 675 581 681
rect 610 675 614 681
rect 648 675 652 681
rect 308 649 312 655
rect 341 649 345 655
rect 374 654 378 660
rect 407 654 411 660
rect 440 654 444 660
rect 478 654 482 660
rect 689 654 693 664
rect 722 654 726 664
rect 755 654 759 664
rect 788 654 792 664
rect 821 654 825 664
rect 519 625 523 635
rect 552 625 556 635
rect 585 625 589 635
rect 618 625 622 635
rect 240 596 285 599
rect 240 595 302 596
rect 316 595 320 609
rect 349 595 353 609
rect 382 604 386 614
rect 415 604 419 614
rect 448 604 452 614
rect 236 584 240 588
rect 272 584 276 595
rect 282 591 309 595
rect 316 591 342 595
rect 349 591 361 595
rect 316 587 320 591
rect 349 587 353 591
rect 185 580 200 584
rect 207 580 240 584
rect -52 441 115 444
rect -52 431 -49 441
rect 8 431 11 441
rect 68 431 71 441
rect 97 435 101 441
rect -58 427 -49 431
rect -128 423 -112 427
rect -44 423 -43 427
rect -128 371 -125 423
rect -61 400 -58 419
rect 7 412 10 419
rect 20 412 23 423
rect 7 409 23 412
rect 69 412 72 419
rect 69 409 83 412
rect 7 406 10 409
rect -52 399 -17 402
rect -121 392 -112 396
rect -105 388 -98 392
rect -105 384 -102 388
rect -52 384 -49 399
rect -105 381 -49 384
rect 7 382 10 394
rect -105 375 -102 381
rect -36 379 10 382
rect -36 375 -33 379
rect 18 372 21 409
rect 69 406 72 409
rect 37 399 45 402
rect 69 382 72 394
rect 26 379 72 382
rect 26 375 29 379
rect -128 367 -113 371
rect -44 367 -43 371
rect 18 368 19 372
rect 79 373 83 409
rect 105 373 109 395
rect 79 369 98 373
rect 105 369 167 373
rect -86 363 -73 367
rect -16 363 -3 367
rect 46 363 59 367
rect 105 365 109 369
rect -76 360 -73 363
rect -6 360 -3 363
rect 56 360 59 363
rect 74 360 85 361
rect -76 357 85 360
rect 81 336 85 357
rect 97 336 101 345
rect 81 333 115 336
rect -53 327 114 330
rect -53 317 -50 327
rect 7 317 10 327
rect 67 317 70 327
rect 96 321 100 327
rect -59 313 -50 317
rect -129 309 -113 313
rect -45 309 -44 313
rect -129 257 -126 309
rect -62 286 -59 305
rect 6 298 9 305
rect 19 298 22 309
rect 6 295 22 298
rect 68 298 71 305
rect 68 295 82 298
rect 6 292 9 295
rect -53 285 -18 288
rect -122 278 -113 282
rect -106 274 -99 278
rect -106 270 -103 274
rect -53 270 -50 285
rect -106 267 -50 270
rect 6 268 9 280
rect -106 261 -103 267
rect -37 265 9 268
rect -37 261 -34 265
rect 17 258 20 295
rect 68 292 71 295
rect 36 285 44 288
rect 68 268 71 280
rect 25 265 71 268
rect 25 261 28 265
rect -129 253 -114 257
rect -45 253 -44 257
rect 17 254 18 258
rect 78 259 82 295
rect 104 259 108 281
rect 78 255 97 259
rect 104 255 156 259
rect -87 249 -74 253
rect -17 249 -4 253
rect 45 249 58 253
rect 104 251 108 255
rect -77 246 -74 249
rect -7 246 -4 249
rect 55 246 58 249
rect 73 246 84 247
rect -77 243 84 246
rect 80 222 84 243
rect 96 222 100 231
rect 80 219 114 222
rect -50 213 117 216
rect -50 203 -47 213
rect 10 203 13 213
rect 70 203 73 213
rect 99 207 103 213
rect -56 199 -47 203
rect -126 195 -110 199
rect -42 195 -41 199
rect -126 143 -123 195
rect -59 172 -56 191
rect 9 184 12 191
rect 22 184 25 195
rect 9 181 25 184
rect 71 184 74 191
rect 71 181 85 184
rect 9 178 12 181
rect -50 171 -15 174
rect -119 164 -110 168
rect -103 160 -96 164
rect -103 156 -100 160
rect -50 156 -47 171
rect -103 153 -47 156
rect 9 154 12 166
rect -103 147 -100 153
rect -34 151 12 154
rect -34 147 -31 151
rect 20 144 23 181
rect 71 178 74 181
rect 39 171 47 174
rect 71 154 74 166
rect 28 151 74 154
rect 28 147 31 151
rect -126 139 -111 143
rect -42 139 -41 143
rect 20 140 21 144
rect 81 145 85 181
rect 107 145 111 167
rect 81 141 100 145
rect 107 141 142 145
rect -84 135 -71 139
rect -14 135 -1 139
rect 48 135 61 139
rect 107 137 111 141
rect -74 132 -71 135
rect -4 132 -1 135
rect 58 132 61 135
rect 76 132 87 133
rect -74 129 87 132
rect 83 108 87 129
rect 99 108 103 117
rect 83 105 117 108
rect -47 99 120 102
rect -47 89 -44 99
rect 13 89 16 99
rect 73 89 76 99
rect 102 93 106 99
rect -53 85 -44 89
rect -123 81 -107 85
rect -39 81 -38 85
rect -123 29 -120 81
rect -56 58 -53 77
rect 12 70 15 77
rect 25 70 28 81
rect 12 67 28 70
rect 74 70 77 77
rect 74 67 88 70
rect 12 64 15 67
rect -47 57 -12 60
rect -116 50 -107 54
rect -100 46 -93 50
rect -100 42 -97 46
rect -47 42 -44 57
rect -100 39 -44 42
rect 12 40 15 52
rect -100 33 -97 39
rect -31 37 15 40
rect -31 33 -28 37
rect 23 30 26 67
rect 74 64 77 67
rect 42 57 50 60
rect 74 40 77 52
rect 31 37 77 40
rect 31 33 34 37
rect -123 25 -108 29
rect -39 25 -38 29
rect 23 26 24 30
rect 84 31 88 67
rect 110 31 114 53
rect 84 27 103 31
rect 110 27 137 31
rect -81 21 -68 25
rect -11 21 2 25
rect 51 21 64 25
rect 110 23 114 27
rect -71 18 -68 21
rect -1 18 2 21
rect 61 18 64 21
rect 79 18 90 19
rect -71 15 90 18
rect 86 -6 90 15
rect 102 -6 106 3
rect 86 -9 120 -6
rect -48 -19 119 -16
rect -48 -29 -45 -19
rect 12 -29 15 -19
rect 72 -29 75 -19
rect 101 -25 105 -19
rect -54 -33 -45 -29
rect -124 -37 -108 -33
rect -40 -37 -39 -33
rect -124 -89 -121 -37
rect -57 -60 -54 -41
rect 11 -48 14 -41
rect 24 -48 27 -37
rect 11 -51 27 -48
rect 73 -48 76 -41
rect 73 -51 87 -48
rect 11 -54 14 -51
rect -48 -61 -13 -58
rect -117 -68 -108 -64
rect -101 -72 -94 -68
rect -101 -76 -98 -72
rect -48 -76 -45 -61
rect -101 -79 -45 -76
rect 11 -78 14 -66
rect -101 -85 -98 -79
rect -32 -81 14 -78
rect -32 -85 -29 -81
rect 22 -88 25 -51
rect 73 -54 76 -51
rect 41 -61 49 -58
rect 73 -78 76 -66
rect 30 -81 76 -78
rect 30 -85 33 -81
rect -124 -93 -109 -89
rect -40 -93 -39 -89
rect 22 -92 23 -88
rect 83 -87 87 -51
rect 109 -87 113 -65
rect 83 -91 102 -87
rect 109 -91 149 -87
rect -82 -97 -69 -93
rect -12 -97 1 -93
rect 50 -97 63 -93
rect 109 -95 113 -91
rect -72 -100 -69 -97
rect -2 -100 1 -97
rect 60 -100 63 -97
rect 78 -100 89 -99
rect -72 -103 89 -100
rect 85 -124 89 -103
rect 101 -124 105 -115
rect 85 -127 119 -124
rect -49 -133 118 -130
rect -49 -143 -46 -133
rect 11 -143 14 -133
rect 71 -143 74 -133
rect 100 -139 104 -133
rect -55 -147 -46 -143
rect -125 -151 -109 -147
rect -41 -151 -40 -147
rect -125 -203 -122 -151
rect -58 -174 -55 -155
rect 10 -162 13 -155
rect 23 -162 26 -151
rect 10 -165 26 -162
rect 72 -162 75 -155
rect 72 -165 86 -162
rect 10 -168 13 -165
rect -49 -175 -14 -172
rect -118 -182 -109 -178
rect -102 -186 -95 -182
rect -102 -190 -99 -186
rect -49 -190 -46 -175
rect -102 -193 -46 -190
rect 10 -192 13 -180
rect -102 -199 -99 -193
rect -33 -195 13 -192
rect -33 -199 -30 -195
rect 21 -202 24 -165
rect 72 -168 75 -165
rect 40 -175 48 -172
rect 72 -192 75 -180
rect 29 -195 75 -192
rect 29 -199 32 -195
rect -125 -207 -110 -203
rect -41 -207 -40 -203
rect 21 -206 22 -202
rect 82 -201 86 -165
rect 108 -201 112 -179
rect 143 -189 149 -91
rect 82 -205 101 -201
rect 108 -205 130 -201
rect -83 -211 -70 -207
rect -13 -211 0 -207
rect 49 -211 62 -207
rect 108 -209 112 -205
rect -73 -214 -70 -211
rect -3 -214 0 -211
rect 59 -214 62 -211
rect 77 -214 88 -213
rect -73 -217 88 -214
rect 84 -238 88 -217
rect 100 -238 104 -229
rect 84 -241 118 -238
rect -46 -247 121 -244
rect -46 -257 -43 -247
rect 14 -257 17 -247
rect 74 -257 77 -247
rect 103 -253 107 -247
rect -52 -261 -43 -257
rect -122 -265 -106 -261
rect -38 -265 -37 -261
rect -122 -317 -119 -265
rect -55 -288 -52 -269
rect 13 -276 16 -269
rect 26 -276 29 -265
rect 13 -279 29 -276
rect 75 -276 78 -269
rect 75 -279 89 -276
rect 13 -282 16 -279
rect -46 -289 -11 -286
rect -115 -296 -106 -292
rect -99 -300 -92 -296
rect -99 -304 -96 -300
rect -46 -304 -43 -289
rect -99 -307 -43 -304
rect 13 -306 16 -294
rect -99 -313 -96 -307
rect -30 -309 16 -306
rect -30 -313 -27 -309
rect 24 -316 27 -279
rect 75 -282 78 -279
rect 43 -289 51 -286
rect 75 -306 78 -294
rect 32 -309 78 -306
rect 32 -313 35 -309
rect -122 -321 -107 -317
rect -38 -321 -37 -317
rect 24 -320 25 -316
rect 85 -315 89 -279
rect 127 -261 130 -205
rect 143 -225 148 -189
rect 143 -231 165 -225
rect 111 -315 115 -293
rect 130 -315 157 -314
rect 85 -319 104 -315
rect 111 -319 158 -315
rect -80 -325 -67 -321
rect -10 -325 3 -321
rect 52 -325 65 -321
rect 111 -323 115 -319
rect 130 -320 158 -319
rect -70 -328 -67 -325
rect 0 -328 3 -325
rect 62 -328 65 -325
rect 80 -328 91 -327
rect -70 -331 91 -328
rect 87 -352 91 -331
rect 103 -352 107 -343
rect 87 -355 121 -352
rect -43 -361 124 -358
rect -43 -371 -40 -361
rect 17 -371 20 -361
rect 77 -371 80 -361
rect 106 -367 110 -361
rect -49 -375 -40 -371
rect -119 -379 -103 -375
rect -35 -379 -34 -375
rect -119 -431 -116 -379
rect -52 -402 -49 -383
rect 16 -390 19 -383
rect 29 -390 32 -379
rect 16 -393 32 -390
rect 78 -390 81 -383
rect 78 -393 92 -390
rect 16 -396 19 -393
rect -43 -403 -8 -400
rect -112 -410 -103 -406
rect -96 -414 -89 -410
rect -96 -418 -93 -414
rect -43 -418 -40 -403
rect -96 -421 -40 -418
rect 16 -420 19 -408
rect -96 -427 -93 -421
rect -27 -423 19 -420
rect -27 -427 -24 -423
rect 27 -430 30 -393
rect 78 -396 81 -393
rect 46 -403 54 -400
rect 78 -420 81 -408
rect 35 -423 81 -420
rect 35 -427 38 -423
rect -119 -435 -104 -431
rect -35 -435 -34 -431
rect 27 -434 28 -430
rect 88 -429 92 -393
rect 154 -379 158 -320
rect 185 -321 188 580
rect 207 576 211 580
rect 199 547 203 556
rect 268 547 272 576
rect 308 547 312 567
rect 341 547 345 567
rect 193 539 360 547
rect 378 537 382 597
rect 401 597 411 601
rect 486 600 490 614
rect 401 556 405 597
rect 444 592 448 597
rect 415 589 448 592
rect 460 596 479 600
rect 486 596 501 600
rect 415 575 421 589
rect 460 578 464 596
rect 486 592 490 596
rect 478 570 482 572
rect 460 559 464 566
rect 401 550 415 556
rect 472 567 482 570
rect 460 540 464 547
rect 284 532 297 536
rect 196 528 257 532
rect 196 446 202 528
rect 280 515 284 524
rect 205 506 229 513
rect 238 512 284 515
rect 244 506 248 512
rect 277 511 284 512
rect 211 500 215 506
rect 219 446 223 460
rect 252 461 256 466
rect 291 461 297 532
rect 378 531 415 537
rect 472 532 476 567
rect 515 539 519 618
rect 548 558 552 618
rect 571 618 581 622
rect 656 621 660 635
rect 571 577 575 618
rect 614 613 618 618
rect 585 610 618 613
rect 630 617 649 621
rect 656 617 671 621
rect 585 596 591 610
rect 630 599 634 617
rect 656 613 660 617
rect 648 591 652 593
rect 630 580 634 587
rect 571 571 585 577
rect 642 588 652 591
rect 630 561 634 568
rect 548 552 585 558
rect 630 542 634 549
rect 515 533 585 539
rect 642 534 646 588
rect 685 549 689 647
rect 718 568 722 647
rect 751 587 755 647
rect 774 647 784 651
rect 859 650 863 664
rect 774 606 778 647
rect 817 642 821 647
rect 788 639 821 642
rect 833 646 852 650
rect 859 646 874 650
rect 788 625 794 639
rect 833 628 837 646
rect 859 642 863 646
rect 851 620 856 622
rect 833 609 837 616
rect 774 600 788 606
rect 846 617 856 620
rect 833 590 837 597
rect 751 581 788 587
rect 833 571 837 578
rect 718 562 788 568
rect 833 552 837 559
rect 685 543 788 549
rect 846 562 850 617
rect 846 558 978 562
rect 846 544 850 558
rect 837 540 850 544
rect 464 528 476 532
rect 634 530 646 534
rect 925 532 947 536
rect 772 527 795 531
rect 521 525 682 527
rect 384 524 682 525
rect 314 522 545 524
rect 314 521 408 522
rect 314 517 371 521
rect 384 518 408 521
rect 417 518 441 522
rect 450 518 474 522
rect 488 518 512 522
rect 521 520 545 522
rect 554 520 578 524
rect 587 520 611 524
rect 620 520 644 524
rect 658 520 682 524
rect 690 523 725 527
rect 320 511 324 517
rect 353 511 357 517
rect 390 512 394 518
rect 423 512 427 518
rect 456 512 460 518
rect 494 512 498 518
rect 527 514 531 520
rect 560 514 564 520
rect 593 514 597 520
rect 626 514 630 520
rect 664 514 668 520
rect 252 458 297 461
rect 252 457 314 458
rect 328 457 332 471
rect 361 457 365 471
rect 398 462 402 472
rect 431 462 435 472
rect 464 462 468 472
rect 248 446 252 450
rect 284 446 288 457
rect 294 453 321 457
rect 328 453 354 457
rect 361 453 373 457
rect 328 449 332 453
rect 361 449 365 453
rect 196 442 212 446
rect 219 442 252 446
rect 196 -186 203 442
rect 219 438 223 442
rect 211 409 215 418
rect 280 409 284 438
rect 320 409 324 429
rect 353 409 357 429
rect 208 402 372 409
rect 337 394 350 398
rect 250 390 310 394
rect 250 308 255 390
rect 333 377 337 386
rect 258 368 282 375
rect 291 374 337 377
rect 297 368 301 374
rect 264 362 268 368
rect 272 308 276 322
rect 305 323 309 328
rect 344 323 350 394
rect 394 395 398 455
rect 417 455 427 459
rect 502 458 506 472
rect 535 464 539 474
rect 568 464 572 474
rect 601 464 605 474
rect 634 464 638 474
rect 417 414 421 455
rect 460 450 464 455
rect 431 447 464 450
rect 476 454 495 458
rect 502 454 517 458
rect 431 433 437 447
rect 476 436 480 454
rect 502 450 506 454
rect 494 428 498 430
rect 476 417 480 424
rect 417 408 431 414
rect 488 425 498 428
rect 476 398 480 405
rect 394 389 431 395
rect 488 390 492 425
rect 480 386 492 390
rect 367 383 424 386
rect 367 379 459 383
rect 373 373 377 379
rect 406 373 410 379
rect 454 364 459 379
rect 531 379 535 457
rect 564 397 568 457
rect 587 457 597 461
rect 672 460 676 474
rect 587 416 591 457
rect 630 452 634 457
rect 601 449 634 452
rect 646 456 665 460
rect 672 456 687 460
rect 601 435 607 449
rect 646 438 650 456
rect 672 452 676 456
rect 664 430 669 432
rect 646 419 650 426
rect 587 410 601 416
rect 659 427 669 430
rect 646 400 650 407
rect 564 391 601 397
rect 646 382 650 388
rect 531 373 601 379
rect 659 374 663 427
rect 690 405 694 523
rect 767 497 772 519
rect 771 493 772 497
rect 711 489 724 493
rect 711 405 715 489
rect 766 462 771 485
rect 790 473 795 527
rect 822 528 878 532
rect 790 466 814 473
rect 796 460 800 466
rect 720 454 724 458
rect 731 444 735 450
rect 723 440 735 444
rect 723 421 727 440
rect 771 425 787 429
rect 723 417 731 421
rect 740 405 744 409
rect 774 405 778 414
rect 782 406 787 425
rect 804 406 808 420
rect 782 402 797 406
rect 804 402 819 406
rect 698 394 699 398
rect 719 394 720 398
rect 748 394 749 398
rect 781 394 782 398
rect 787 394 791 402
rect 804 398 808 402
rect 687 374 691 378
rect 708 374 712 378
rect 737 374 741 378
rect 770 374 774 378
rect 797 374 801 378
rect 650 371 801 374
rect 822 377 826 528
rect 920 503 925 524
rect 924 499 925 503
rect 842 495 877 499
rect 842 377 846 495
rect 919 469 924 491
rect 923 465 924 469
rect 863 461 876 465
rect 863 377 867 461
rect 918 434 923 457
rect 942 445 947 532
rect 942 438 966 445
rect 948 432 952 438
rect 872 426 876 430
rect 883 416 887 422
rect 875 412 887 416
rect 875 393 879 412
rect 923 397 939 401
rect 875 389 883 393
rect 892 377 896 379
rect 926 377 930 386
rect 934 378 939 397
rect 956 378 960 392
rect 934 374 949 378
rect 956 374 971 378
rect 650 370 663 371
rect 440 361 694 364
rect 440 357 464 361
rect 473 357 497 361
rect 506 357 530 361
rect 544 357 568 361
rect 305 320 350 323
rect 305 319 367 320
rect 381 319 385 333
rect 414 319 418 333
rect 446 351 450 357
rect 479 351 483 357
rect 512 351 516 357
rect 550 351 554 357
rect 657 354 681 358
rect 301 308 305 312
rect 337 308 341 319
rect 347 315 374 319
rect 381 315 407 319
rect 414 315 426 319
rect 381 311 385 315
rect 414 311 418 315
rect 209 304 265 308
rect 272 304 305 308
rect 209 -53 216 304
rect 272 300 276 304
rect 265 271 269 280
rect 334 271 338 300
rect 454 301 458 311
rect 487 301 491 311
rect 520 301 524 311
rect 374 271 378 291
rect 407 271 411 291
rect 227 266 425 271
rect 227 263 441 266
rect 337 256 350 260
rect 250 252 310 256
rect 250 170 255 252
rect 333 239 337 248
rect 258 230 282 237
rect 291 236 337 239
rect 297 230 301 236
rect 264 224 268 230
rect 272 170 276 184
rect 305 185 309 190
rect 344 185 350 256
rect 367 241 430 248
rect 373 235 377 241
rect 406 235 410 241
rect 305 182 350 185
rect 305 181 367 182
rect 381 181 385 195
rect 414 181 418 195
rect 427 195 430 241
rect 435 221 441 263
rect 450 234 454 294
rect 473 294 483 298
rect 558 297 562 311
rect 597 350 610 354
rect 473 253 477 294
rect 516 289 520 294
rect 487 286 520 289
rect 532 293 551 297
rect 558 293 573 297
rect 487 272 493 286
rect 532 275 536 293
rect 558 289 562 293
rect 550 267 555 269
rect 532 256 536 263
rect 473 247 487 253
rect 545 264 555 267
rect 597 266 601 350
rect 652 323 657 346
rect 676 334 681 354
rect 691 334 694 361
rect 796 346 801 371
rect 830 366 831 370
rect 850 366 851 370
rect 871 366 872 370
rect 900 366 901 370
rect 933 366 934 370
rect 939 366 943 374
rect 956 370 960 374
rect 819 346 823 350
rect 839 346 843 350
rect 860 346 864 350
rect 889 346 893 350
rect 922 346 926 350
rect 949 346 953 350
rect 975 346 978 558
rect 1091 472 1258 475
rect 1091 462 1094 472
rect 1151 462 1154 472
rect 1211 462 1214 472
rect 1240 466 1244 472
rect 1085 458 1094 462
rect 1015 454 1031 458
rect 1099 454 1100 458
rect 1015 402 1018 454
rect 1082 431 1085 450
rect 1150 443 1153 450
rect 1163 443 1166 454
rect 1150 440 1166 443
rect 1212 443 1215 450
rect 1212 440 1226 443
rect 1150 437 1153 440
rect 1091 430 1126 433
rect 1022 423 1031 427
rect 1038 419 1045 423
rect 1038 415 1041 419
rect 1091 415 1094 430
rect 1038 412 1094 415
rect 1150 413 1153 425
rect 1038 406 1041 412
rect 1107 410 1153 413
rect 1107 406 1110 410
rect 1161 403 1164 440
rect 1212 437 1215 440
rect 1180 430 1188 433
rect 1212 413 1215 425
rect 1169 410 1215 413
rect 1169 406 1172 410
rect 1015 398 1030 402
rect 1099 398 1100 402
rect 1161 399 1162 403
rect 1222 404 1226 440
rect 1248 404 1252 426
rect 1222 400 1241 404
rect 1248 400 1258 404
rect 1015 376 1018 398
rect 1057 394 1070 398
rect 1127 394 1140 398
rect 1189 394 1202 398
rect 1248 396 1252 400
rect 1067 391 1070 394
rect 1137 391 1140 394
rect 1199 391 1202 394
rect 1217 391 1228 392
rect 1067 388 1228 391
rect 1224 367 1228 388
rect 1240 367 1244 376
rect 1224 364 1258 367
rect 796 343 978 346
rect 717 337 807 340
rect 676 327 700 334
rect 682 321 686 327
rect 607 315 610 319
rect 617 305 621 311
rect 609 301 621 305
rect 609 282 613 301
rect 657 286 673 290
rect 609 278 617 282
rect 532 237 536 244
rect 450 228 487 234
rect 545 229 549 264
rect 626 266 630 269
rect 660 266 664 275
rect 668 267 673 286
rect 690 267 694 281
rect 668 263 683 267
rect 690 263 705 267
rect 605 255 606 259
rect 634 255 635 259
rect 667 255 668 259
rect 673 255 677 263
rect 690 259 694 263
rect 717 262 722 337
rect 768 329 772 337
rect 725 322 749 329
rect 803 326 807 337
rect 834 333 891 340
rect 840 327 844 333
rect 873 327 877 333
rect 731 316 735 322
rect 739 262 743 276
rect 717 258 732 262
rect 739 258 754 262
rect 739 254 743 258
rect 594 235 598 239
rect 623 235 627 239
rect 656 235 660 239
rect 683 235 687 239
rect 594 232 687 235
rect 749 248 754 258
rect 764 261 768 282
rect 815 286 833 290
rect 772 273 776 282
rect 806 276 812 278
rect 829 273 833 286
rect 848 273 852 287
rect 881 273 885 287
rect 772 269 841 273
rect 848 269 874 273
rect 881 269 896 273
rect 804 261 807 269
rect 764 257 772 261
rect 810 258 819 261
rect 784 248 788 253
rect 810 248 813 258
rect 749 245 813 248
rect 749 244 788 245
rect 536 228 549 229
rect 683 228 688 232
rect 536 225 688 228
rect 732 225 736 234
rect 812 233 816 240
rect 831 250 835 269
rect 848 265 852 269
rect 881 265 885 269
rect 828 247 835 250
rect 892 253 896 269
rect 841 225 845 245
rect 874 225 878 245
rect 902 225 910 343
rect 544 221 549 225
rect 435 218 549 221
rect 683 219 688 225
rect 726 219 910 225
rect 683 217 910 219
rect 683 214 732 217
rect 480 195 700 196
rect 427 192 700 195
rect 480 191 700 192
rect 480 185 485 191
rect 504 189 700 191
rect 510 183 514 189
rect 301 170 305 174
rect 337 170 341 181
rect 347 177 374 181
rect 381 177 407 181
rect 414 177 438 181
rect 381 173 385 177
rect 414 173 418 177
rect 238 166 265 170
rect 272 166 305 170
rect 238 81 243 166
rect 272 162 276 166
rect 264 133 268 142
rect 333 133 337 162
rect 373 133 377 153
rect 406 133 410 153
rect 257 125 424 133
rect 272 105 276 125
rect 305 105 309 125
rect 314 100 321 103
rect 264 81 268 85
rect 297 81 301 85
rect 314 81 318 100
rect 414 116 418 125
rect 361 105 400 106
rect 336 102 400 105
rect 336 92 339 102
rect 361 97 365 102
rect 330 89 339 92
rect 377 89 385 93
rect 342 81 345 89
rect 238 77 268 81
rect 275 77 301 81
rect 308 77 377 81
rect 264 63 268 77
rect 297 63 301 77
rect 316 64 320 77
rect 337 72 343 74
rect 373 68 377 77
rect 316 60 334 64
rect 381 68 385 89
rect 395 92 400 102
rect 421 98 424 125
rect 427 128 431 177
rect 445 167 449 173
rect 437 163 449 167
rect 437 144 441 163
rect 485 148 501 152
rect 437 140 445 144
rect 488 128 492 137
rect 427 124 454 128
rect 496 129 501 148
rect 518 129 522 143
rect 630 139 643 143
rect 543 135 603 139
rect 496 125 511 129
rect 518 125 533 129
rect 462 117 463 121
rect 495 117 496 121
rect 501 117 505 125
rect 518 121 522 125
rect 421 97 438 98
rect 450 97 454 101
rect 483 97 487 101
rect 510 98 514 101
rect 510 97 531 98
rect 406 92 410 96
rect 421 95 531 97
rect 435 94 514 95
rect 395 88 410 92
rect 417 88 432 92
rect 406 74 410 88
rect 414 28 418 34
rect 427 38 432 88
rect 427 30 505 38
rect 272 17 276 23
rect 305 17 309 23
rect 258 10 315 17
rect 342 6 346 24
rect 400 21 424 28
rect 377 6 381 21
rect 427 6 432 30
rect 470 25 505 30
rect 470 9 505 22
rect 527 9 531 95
rect 543 53 548 135
rect 626 122 630 131
rect 551 113 575 120
rect 584 119 630 122
rect 590 113 594 119
rect 557 107 561 113
rect 565 53 569 67
rect 598 68 602 73
rect 637 68 643 139
rect 692 131 700 189
rect 660 124 717 131
rect 666 118 670 124
rect 699 118 703 124
rect 598 65 643 68
rect 598 64 660 65
rect 674 64 678 78
rect 707 64 711 78
rect 594 53 598 57
rect 630 53 634 64
rect 640 60 667 64
rect 674 60 700 64
rect 707 60 719 64
rect 674 56 678 60
rect 707 56 711 60
rect 743 58 762 66
rect 543 49 558 53
rect 565 49 598 53
rect 565 45 569 49
rect 557 16 561 25
rect 626 16 630 45
rect 666 16 670 36
rect 699 16 703 36
rect 551 13 718 16
rect 551 12 726 13
rect 551 9 727 12
rect 342 2 432 6
rect 527 8 727 9
rect 527 5 558 8
rect 533 -1 537 5
rect 627 1 640 5
rect 257 -4 537 -1
rect 257 -9 424 -4
rect 533 -5 537 -4
rect 540 -3 600 1
rect 272 -29 276 -9
rect 305 -29 309 -9
rect 314 -34 321 -31
rect 264 -53 268 -49
rect 297 -53 301 -49
rect 314 -53 318 -34
rect 414 -18 418 -9
rect 361 -29 400 -28
rect 336 -32 400 -29
rect 336 -42 339 -32
rect 361 -37 365 -32
rect 330 -45 339 -42
rect 377 -45 385 -41
rect 342 -53 345 -45
rect 209 -57 268 -53
rect 275 -57 301 -53
rect 308 -57 377 -53
rect 264 -71 268 -57
rect 297 -71 301 -57
rect 316 -70 320 -57
rect 337 -62 343 -60
rect 373 -66 377 -57
rect 316 -74 334 -70
rect 381 -66 385 -45
rect 395 -42 400 -32
rect 406 -42 410 -38
rect 395 -46 410 -42
rect 417 -46 432 -42
rect 406 -60 410 -46
rect 414 -106 418 -100
rect 427 -101 432 -46
rect 540 -85 545 -3
rect 623 -16 627 -7
rect 548 -25 572 -18
rect 581 -19 627 -16
rect 587 -25 591 -19
rect 554 -31 558 -25
rect 562 -85 566 -71
rect 595 -70 599 -65
rect 634 -70 640 1
rect 657 -14 714 -7
rect 663 -20 667 -14
rect 696 -20 700 -14
rect 595 -73 640 -70
rect 595 -74 657 -73
rect 671 -74 675 -60
rect 704 -74 708 -60
rect 591 -85 595 -81
rect 627 -85 631 -74
rect 637 -78 664 -74
rect 671 -78 697 -74
rect 704 -78 716 -74
rect 671 -82 675 -78
rect 704 -82 708 -78
rect 540 -89 555 -85
rect 562 -89 595 -85
rect 562 -93 566 -89
rect 470 -101 505 -99
rect 272 -117 276 -111
rect 305 -117 309 -111
rect 258 -124 315 -117
rect 342 -128 346 -110
rect 400 -113 424 -106
rect 427 -107 505 -101
rect 377 -128 381 -113
rect 427 -128 432 -107
rect 470 -112 505 -107
rect 470 -127 505 -115
rect 554 -122 558 -113
rect 623 -122 627 -93
rect 663 -122 667 -102
rect 696 -122 700 -102
rect 548 -125 715 -122
rect 724 -125 727 8
rect 777 -3 867 1
rect 744 -80 756 -72
rect 777 -85 782 -3
rect 828 -18 832 -3
rect 789 -25 813 -18
rect 863 -21 867 -3
rect 791 -31 795 -25
rect 799 -85 803 -71
rect 777 -89 792 -85
rect 799 -89 814 -85
rect 799 -93 803 -89
rect 809 -99 814 -89
rect 824 -86 828 -65
rect 875 -61 893 -57
rect 832 -74 836 -65
rect 866 -71 872 -69
rect 889 -74 893 -61
rect 832 -78 894 -74
rect 864 -86 867 -78
rect 824 -90 832 -86
rect 870 -89 879 -86
rect 844 -99 848 -94
rect 870 -99 873 -89
rect 809 -102 873 -99
rect 809 -103 848 -102
rect 792 -122 796 -113
rect 872 -114 876 -109
rect 891 -97 894 -78
rect 888 -100 894 -97
rect 903 -122 910 217
rect 1072 152 1239 155
rect 1072 142 1075 152
rect 1132 142 1135 152
rect 1192 142 1195 152
rect 1221 146 1225 152
rect 1066 138 1075 142
rect 996 134 1012 138
rect 1080 134 1081 138
rect 996 82 999 134
rect 1063 111 1066 130
rect 1131 123 1134 130
rect 1144 123 1147 134
rect 1131 120 1147 123
rect 1193 123 1196 130
rect 1193 120 1207 123
rect 1131 117 1134 120
rect 1072 110 1107 113
rect 1003 103 1012 107
rect 1019 99 1026 103
rect 1019 95 1022 99
rect 1072 95 1075 110
rect 1019 92 1075 95
rect 1131 93 1134 105
rect 1019 86 1022 92
rect 1088 90 1134 93
rect 1088 86 1091 90
rect 1142 83 1145 120
rect 1193 117 1196 120
rect 1161 110 1169 113
rect 1193 93 1196 105
rect 1150 90 1196 93
rect 1150 86 1153 90
rect 996 78 1011 82
rect 1080 78 1081 82
rect 1142 79 1143 83
rect 1203 84 1207 120
rect 1229 84 1233 106
rect 1203 80 1222 84
rect 1229 80 1239 84
rect 1038 74 1051 78
rect 1108 74 1121 78
rect 1170 74 1183 78
rect 1229 76 1233 80
rect 1048 71 1051 74
rect 1118 71 1121 74
rect 1180 71 1183 74
rect 1198 71 1209 72
rect 1048 68 1209 71
rect 1205 47 1209 68
rect 1221 47 1225 56
rect 1205 44 1239 47
rect 1071 38 1238 41
rect 1071 28 1074 38
rect 1131 28 1134 38
rect 1191 28 1194 38
rect 1220 32 1224 38
rect 1065 24 1074 28
rect 995 20 1011 24
rect 1079 20 1080 24
rect 995 -32 998 20
rect 1062 -3 1065 16
rect 1130 9 1133 16
rect 1143 9 1146 20
rect 1130 6 1146 9
rect 1192 9 1195 16
rect 1192 6 1206 9
rect 1130 3 1133 6
rect 1071 -4 1106 -1
rect 1002 -11 1011 -7
rect 1018 -15 1025 -11
rect 1018 -19 1021 -15
rect 1071 -19 1074 -4
rect 1018 -22 1074 -19
rect 1130 -21 1133 -9
rect 1018 -28 1021 -22
rect 1087 -24 1133 -21
rect 1087 -28 1090 -24
rect 1141 -31 1144 6
rect 1192 3 1195 6
rect 1160 -4 1168 -1
rect 1192 -21 1195 -9
rect 1149 -24 1195 -21
rect 1149 -28 1152 -24
rect 995 -36 1010 -32
rect 1079 -36 1080 -32
rect 1141 -35 1142 -31
rect 1202 -30 1206 6
rect 1228 -30 1232 -8
rect 1202 -34 1221 -30
rect 1228 -34 1238 -30
rect 1037 -40 1050 -36
rect 1107 -40 1120 -36
rect 1169 -40 1182 -36
rect 1228 -38 1232 -34
rect 1047 -43 1050 -40
rect 1117 -43 1120 -40
rect 1179 -43 1182 -40
rect 1197 -43 1208 -42
rect 1047 -46 1208 -43
rect 1204 -67 1208 -46
rect 1220 -67 1224 -58
rect 1204 -70 1238 -67
rect 1074 -76 1241 -73
rect 1074 -86 1077 -76
rect 1134 -86 1137 -76
rect 1194 -86 1197 -76
rect 1223 -82 1227 -76
rect 1068 -90 1077 -86
rect 342 -132 432 -128
rect 523 -129 727 -125
rect 317 -136 425 -135
rect 523 -136 530 -129
rect 548 -130 727 -129
rect 786 -129 910 -122
rect 998 -94 1014 -90
rect 1082 -94 1083 -90
rect 786 -130 904 -129
rect 317 -143 530 -136
rect 630 -137 643 -133
rect 543 -141 603 -137
rect 315 -168 322 -165
rect 315 -186 319 -168
rect 415 -152 419 -143
rect 362 -163 401 -162
rect 337 -166 401 -163
rect 337 -176 340 -166
rect 362 -171 366 -166
rect 331 -179 340 -176
rect 378 -179 386 -175
rect 196 -187 319 -186
rect 343 -187 346 -179
rect 196 -191 378 -187
rect 317 -204 321 -191
rect 338 -196 344 -194
rect 374 -200 378 -191
rect 317 -208 335 -204
rect 382 -200 386 -179
rect 396 -176 401 -166
rect 407 -176 411 -172
rect 396 -180 411 -176
rect 418 -180 433 -176
rect 407 -194 411 -180
rect 415 -240 419 -234
rect 428 -240 433 -180
rect 543 -223 548 -141
rect 626 -154 630 -145
rect 551 -163 575 -156
rect 584 -157 630 -154
rect 590 -163 594 -157
rect 557 -169 561 -163
rect 565 -223 569 -209
rect 598 -208 602 -203
rect 637 -208 643 -137
rect 598 -211 643 -208
rect 774 -137 864 -133
rect 998 -135 1001 -94
rect 1065 -117 1068 -98
rect 1133 -105 1136 -98
rect 1146 -105 1149 -94
rect 1133 -108 1149 -105
rect 1195 -105 1198 -98
rect 1195 -108 1209 -105
rect 1133 -111 1136 -108
rect 1074 -118 1109 -115
rect 1005 -125 1014 -121
rect 774 -211 779 -137
rect 825 -152 829 -137
rect 782 -159 806 -152
rect 860 -155 864 -137
rect 968 -138 1001 -135
rect 788 -165 792 -159
rect 598 -212 766 -211
rect 594 -223 598 -219
rect 630 -223 634 -212
rect 640 -216 766 -212
rect 660 -217 766 -216
rect 746 -219 766 -217
rect 771 -219 779 -211
rect 796 -219 800 -205
rect 774 -223 789 -219
rect 796 -223 811 -219
rect 543 -227 558 -223
rect 565 -227 598 -223
rect 796 -227 800 -223
rect 565 -231 569 -227
rect 470 -240 505 -237
rect 343 -262 347 -244
rect 401 -247 425 -240
rect 428 -246 505 -240
rect 378 -262 382 -247
rect 428 -262 433 -246
rect 470 -249 505 -246
rect 343 -266 433 -262
rect 470 -265 505 -252
rect 557 -260 561 -251
rect 626 -260 630 -231
rect 806 -233 811 -223
rect 821 -220 825 -199
rect 872 -195 890 -191
rect 829 -208 833 -199
rect 863 -205 869 -203
rect 886 -205 890 -195
rect 968 -205 973 -138
rect 998 -146 1001 -138
rect 1021 -129 1028 -125
rect 1021 -133 1024 -129
rect 1074 -133 1077 -118
rect 1021 -136 1077 -133
rect 1133 -135 1136 -123
rect 1021 -142 1024 -136
rect 1090 -138 1136 -135
rect 1090 -142 1093 -138
rect 1144 -145 1147 -108
rect 1195 -111 1198 -108
rect 1163 -118 1171 -115
rect 1195 -135 1198 -123
rect 1152 -138 1198 -135
rect 1152 -142 1155 -138
rect 998 -150 1013 -146
rect 1082 -150 1083 -146
rect 1144 -149 1145 -145
rect 1205 -144 1209 -108
rect 1231 -144 1235 -122
rect 1205 -148 1224 -144
rect 1231 -148 1241 -144
rect 1040 -154 1053 -150
rect 1110 -154 1123 -150
rect 1172 -154 1185 -150
rect 1231 -152 1235 -148
rect 1050 -157 1053 -154
rect 1120 -157 1123 -154
rect 1182 -157 1185 -154
rect 1200 -157 1211 -156
rect 1050 -160 1211 -157
rect 1207 -181 1211 -160
rect 1223 -181 1227 -172
rect 1207 -184 1241 -181
rect 1077 -190 1244 -187
rect 1077 -200 1080 -190
rect 1137 -200 1140 -190
rect 1197 -200 1200 -190
rect 1226 -196 1230 -190
rect 1071 -204 1080 -200
rect 886 -208 973 -205
rect 829 -210 973 -208
rect 1001 -208 1017 -204
rect 1085 -208 1086 -204
rect 829 -212 891 -210
rect 861 -220 864 -212
rect 821 -224 829 -220
rect 867 -223 876 -220
rect 841 -233 845 -228
rect 867 -233 870 -223
rect 806 -236 870 -233
rect 806 -237 845 -236
rect 788 -256 792 -247
rect 869 -248 873 -243
rect 888 -231 891 -212
rect 885 -234 891 -231
rect 551 -268 660 -260
rect 782 -264 891 -256
rect 1001 -260 1004 -208
rect 1068 -231 1071 -212
rect 1136 -219 1139 -212
rect 1149 -219 1152 -208
rect 1136 -222 1152 -219
rect 1198 -219 1201 -212
rect 1198 -222 1212 -219
rect 1136 -225 1139 -222
rect 1077 -232 1112 -229
rect 1008 -239 1017 -235
rect 1024 -243 1031 -239
rect 1024 -247 1027 -243
rect 1077 -247 1080 -232
rect 1024 -250 1080 -247
rect 1136 -249 1139 -237
rect 1024 -256 1027 -250
rect 1093 -252 1139 -249
rect 1093 -256 1096 -252
rect 1147 -259 1150 -222
rect 1198 -225 1201 -222
rect 1166 -232 1174 -229
rect 1198 -249 1201 -237
rect 1155 -252 1201 -249
rect 1155 -256 1158 -252
rect 1001 -264 1016 -260
rect 1085 -264 1086 -260
rect 1147 -263 1148 -259
rect 1208 -258 1212 -222
rect 1234 -258 1238 -236
rect 1208 -262 1227 -258
rect 1234 -262 1244 -258
rect 317 -277 425 -269
rect 787 -271 911 -267
rect 630 -275 643 -271
rect 315 -302 322 -299
rect 315 -321 319 -302
rect 415 -286 419 -277
rect 362 -297 401 -296
rect 337 -300 401 -297
rect 337 -310 340 -300
rect 362 -305 366 -300
rect 331 -313 340 -310
rect 378 -313 386 -309
rect 343 -321 346 -313
rect 185 -325 378 -321
rect 256 -326 322 -325
rect 317 -338 321 -326
rect 338 -330 344 -328
rect 374 -334 378 -325
rect 317 -342 335 -338
rect 154 -387 175 -379
rect 114 -429 118 -407
rect 317 -425 320 -342
rect 382 -334 386 -313
rect 396 -310 401 -300
rect 543 -279 603 -275
rect 407 -310 411 -306
rect 396 -314 411 -310
rect 418 -314 433 -310
rect 407 -328 411 -314
rect 415 -374 419 -368
rect 343 -396 347 -378
rect 401 -381 425 -374
rect 378 -396 382 -381
rect 428 -382 433 -314
rect 543 -361 548 -279
rect 626 -292 630 -283
rect 551 -301 575 -294
rect 584 -295 630 -292
rect 590 -301 594 -295
rect 557 -307 561 -301
rect 565 -361 569 -347
rect 598 -346 602 -341
rect 637 -346 643 -275
rect 660 -290 717 -283
rect 666 -296 670 -290
rect 699 -296 703 -290
rect 598 -349 643 -346
rect 598 -350 660 -349
rect 674 -350 678 -336
rect 707 -350 711 -336
rect 594 -361 598 -357
rect 630 -361 634 -350
rect 640 -354 667 -350
rect 674 -354 700 -350
rect 707 -354 719 -350
rect 674 -358 678 -354
rect 707 -358 711 -354
rect 746 -356 774 -348
rect 787 -353 792 -271
rect 838 -286 842 -271
rect 795 -293 819 -286
rect 873 -289 877 -271
rect 801 -299 805 -293
rect 809 -353 813 -339
rect 543 -365 558 -361
rect 565 -365 598 -361
rect 565 -369 569 -365
rect 470 -382 505 -377
rect 428 -388 505 -382
rect 428 -396 433 -388
rect 470 -390 505 -388
rect 343 -400 433 -396
rect 470 -406 505 -393
rect 557 -398 561 -389
rect 626 -398 630 -369
rect 787 -357 802 -353
rect 809 -357 824 -353
rect 666 -398 670 -378
rect 699 -398 703 -378
rect 551 -406 718 -398
rect 787 -404 791 -357
rect 809 -361 813 -357
rect 819 -367 824 -357
rect 834 -354 838 -333
rect 885 -329 903 -325
rect 842 -342 846 -333
rect 876 -339 882 -337
rect 899 -342 903 -329
rect 1011 -342 1015 -264
rect 1043 -268 1056 -264
rect 1113 -268 1126 -264
rect 1175 -268 1188 -264
rect 1234 -266 1238 -262
rect 1053 -271 1056 -268
rect 1123 -271 1126 -268
rect 1185 -271 1188 -268
rect 1203 -271 1214 -270
rect 1053 -274 1214 -271
rect 842 -346 1015 -342
rect 874 -354 877 -346
rect 834 -358 842 -354
rect 880 -357 889 -354
rect 854 -367 858 -362
rect 880 -367 883 -357
rect 819 -370 883 -367
rect 819 -371 858 -370
rect 801 -390 805 -381
rect 883 -382 886 -377
rect 901 -365 905 -346
rect 898 -368 905 -365
rect 795 -392 905 -390
rect 1186 -392 1195 -274
rect 1210 -295 1214 -274
rect 1226 -295 1230 -286
rect 1210 -298 1244 -295
rect 795 -396 1195 -392
rect 795 -397 1192 -396
rect 795 -398 905 -397
rect 787 -414 794 -404
rect 790 -425 794 -414
rect 317 -428 794 -425
rect 88 -433 107 -429
rect 114 -433 189 -429
rect -77 -439 -64 -435
rect -7 -439 6 -435
rect 55 -439 68 -435
rect 114 -437 118 -433
rect -67 -442 -64 -439
rect 3 -442 6 -439
rect 65 -442 68 -439
rect 83 -442 94 -441
rect -67 -445 94 -442
rect 90 -466 94 -445
rect 106 -466 110 -457
rect 321 -466 554 -465
rect 90 -468 554 -466
rect 90 -469 324 -468
<< metal2 >>
rect 208 655 302 662
rect 208 651 216 655
rect 694 654 722 659
rect 727 654 755 659
rect 760 654 788 659
rect 793 654 821 659
rect 826 654 842 659
rect 838 651 842 654
rect 872 645 931 650
rect 265 607 272 644
rect 524 625 552 630
rect 557 625 585 630
rect 590 625 618 630
rect 623 625 639 630
rect 635 622 639 625
rect 665 617 898 623
rect 172 603 272 607
rect 387 604 415 609
rect 420 604 448 609
rect 453 604 469 609
rect -47 397 -42 426
rect -116 395 -42 397
rect 40 395 43 402
rect -116 392 45 395
rect -47 391 45 392
rect -47 371 -42 391
rect -48 283 -43 312
rect -117 281 -43 283
rect 39 281 42 288
rect -117 278 44 281
rect -48 277 44 278
rect -48 257 -43 277
rect -45 169 -40 198
rect -114 167 -40 169
rect 42 167 45 174
rect -114 164 47 167
rect -45 163 47 164
rect -45 143 -40 163
rect -42 55 -37 84
rect -111 53 -37 55
rect 45 53 48 60
rect -111 50 50 53
rect -42 49 50 50
rect -42 29 -37 49
rect -43 -63 -38 -34
rect -112 -65 -38 -63
rect 44 -65 47 -58
rect -112 -68 49 -65
rect -43 -69 49 -68
rect -43 -89 -38 -69
rect -44 -177 -39 -148
rect -113 -179 -39 -177
rect 43 -179 46 -172
rect -113 -182 48 -179
rect -44 -183 48 -182
rect -44 -203 -39 -183
rect -41 -291 -36 -262
rect 172 -267 177 603
rect 465 601 469 604
rect 358 590 364 597
rect 498 596 873 601
rect 358 585 851 590
rect 842 583 851 585
rect 527 567 692 568
rect 185 561 692 567
rect 249 550 405 556
rect 249 528 255 550
rect 220 517 314 524
rect 220 513 228 517
rect 277 500 410 505
rect 277 483 284 500
rect 842 494 850 583
rect 181 477 284 483
rect 181 -128 192 477
rect 403 462 431 467
rect 436 462 464 467
rect 469 462 485 467
rect 540 464 568 469
rect 573 464 601 469
rect 606 464 634 469
rect 639 464 655 469
rect 481 459 485 462
rect 651 461 655 464
rect 867 460 873 596
rect 682 453 719 458
rect 417 443 568 448
rect 417 415 422 443
rect 198 410 399 415
rect 415 397 423 415
rect 303 390 423 397
rect 273 379 367 386
rect 273 375 281 379
rect 431 373 437 439
rect 715 409 719 453
rect 893 448 898 617
rect 867 445 898 448
rect 715 405 740 409
rect 699 394 715 398
rect 720 394 744 398
rect 749 394 777 398
rect 782 394 787 398
rect 671 373 677 391
rect 867 381 871 445
rect 867 377 892 381
rect 926 379 931 645
rect 1096 428 1101 457
rect 1027 426 1101 428
rect 1183 426 1186 433
rect 1027 423 1188 426
rect 1096 422 1188 423
rect 1096 402 1101 422
rect 965 374 1017 380
rect 337 368 681 373
rect 459 301 487 306
rect 492 301 520 306
rect 525 301 541 306
rect 537 298 541 301
rect 273 241 367 248
rect 273 237 281 241
rect 572 165 576 368
rect 831 366 846 370
rect 851 366 867 370
rect 872 366 896 370
rect 901 366 929 370
rect 934 366 939 370
rect 597 333 710 338
rect 601 270 605 319
rect 601 266 626 270
rect 606 255 630 259
rect 635 255 663 259
rect 668 255 673 259
rect 705 212 710 333
rect 740 333 834 340
rect 740 329 748 333
rect 806 271 812 276
rect 769 265 812 271
rect 807 232 812 265
rect 705 208 773 212
rect 488 160 733 165
rect 488 135 492 160
rect 566 126 660 131
rect 337 85 342 118
rect 463 117 491 121
rect 496 117 501 121
rect 566 120 574 126
rect 337 79 381 85
rect 386 79 463 85
rect 337 73 343 79
rect 455 21 463 79
rect 615 21 620 114
rect 727 66 733 160
rect 720 58 740 66
rect 768 21 773 208
rect 1077 108 1082 137
rect 1008 106 1082 108
rect 1164 106 1167 113
rect 1008 103 1169 106
rect 1077 102 1169 103
rect 1077 82 1082 102
rect 401 17 409 21
rect 315 10 409 17
rect 455 14 494 21
rect 502 16 620 21
rect 728 16 773 21
rect 563 -12 657 -7
rect 337 -49 342 -16
rect 563 -18 571 -12
rect 337 -55 381 -49
rect 386 -55 452 -49
rect 337 -60 343 -55
rect 401 -117 409 -113
rect 315 -124 409 -117
rect 443 -116 452 -55
rect 610 -116 617 -23
rect 728 -72 736 16
rect 1076 -6 1081 23
rect 1007 -8 1081 -6
rect 1163 -8 1166 -1
rect 1007 -11 1168 -8
rect 1076 -12 1168 -11
rect 1076 -32 1081 -12
rect 720 -80 741 -72
rect 866 -76 872 -71
rect 443 -123 491 -116
rect 501 -121 617 -116
rect 728 -128 735 -80
rect 829 -82 872 -76
rect 867 -115 872 -82
rect 1079 -120 1084 -91
rect 1010 -122 1084 -120
rect 1166 -122 1169 -115
rect 1010 -125 1171 -122
rect 181 -135 735 -128
rect 1079 -126 1171 -125
rect 1079 -146 1084 -126
rect 338 -183 343 -150
rect 338 -189 382 -183
rect 387 -189 451 -183
rect 338 -194 344 -189
rect 444 -254 451 -189
rect 619 -254 624 -161
rect 863 -210 869 -205
rect 723 -219 743 -211
rect 826 -216 869 -210
rect 444 -259 496 -254
rect 503 -259 624 -254
rect 731 -267 739 -219
rect 864 -249 869 -216
rect 1082 -234 1087 -205
rect 1013 -236 1087 -234
rect 1169 -236 1172 -229
rect 1013 -239 1174 -236
rect 1082 -240 1174 -239
rect 1082 -260 1087 -240
rect 172 -268 660 -267
rect 719 -268 739 -267
rect 172 -272 739 -268
rect -110 -293 -36 -291
rect 46 -293 49 -286
rect -110 -296 51 -293
rect -41 -297 51 -296
rect -41 -317 -36 -297
rect 338 -317 343 -284
rect 566 -287 660 -283
rect 566 -294 574 -287
rect 338 -323 382 -317
rect 387 -323 450 -317
rect 338 -328 344 -323
rect -38 -405 -33 -376
rect 442 -394 450 -323
rect 617 -393 622 -299
rect 876 -344 882 -339
rect 723 -356 743 -348
rect 839 -350 882 -344
rect 877 -383 882 -350
rect 442 -400 496 -394
rect 503 -397 622 -393
rect -107 -407 -33 -405
rect 49 -407 52 -400
rect -107 -410 54 -407
rect -38 -411 54 -410
rect -38 -431 -33 -411
<< metal3 >>
rect 574 572 756 579
rect 401 550 554 556
rect 370 453 453 458
rect -117 283 -112 397
rect -117 278 -109 283
rect -114 169 -109 278
rect -114 164 -107 169
rect -112 53 -107 164
rect 78 104 85 447
rect 448 441 453 453
rect 574 445 579 572
rect 1204 472 1212 478
rect 810 467 1212 472
rect 810 466 961 467
rect 636 449 642 459
rect 448 437 556 441
rect 563 440 580 445
rect 636 444 714 449
rect 551 430 556 437
rect 394 421 534 426
rect 551 425 778 430
rect 394 410 399 421
rect 774 406 778 425
rect 78 98 87 104
rect -112 50 -106 53
rect -111 -63 -106 50
rect -112 -66 -106 -63
rect 82 -13 87 98
rect 111 -2 117 340
rect 111 -9 119 -2
rect -112 -177 -107 -66
rect -112 -182 -105 -177
rect -110 -291 -105 -182
rect -110 -296 -102 -291
rect -107 -410 -102 -296
rect 82 -362 89 -13
rect 114 -120 119 -9
rect 114 -127 121 -120
rect -107 -471 -103 -410
rect 115 -467 121 -127
rect 131 -141 136 33
rect 144 -92 148 148
rect 154 -5 159 264
rect 166 45 171 371
rect 834 337 840 466
rect 954 441 961 466
rect 425 315 609 320
rect 566 293 665 298
rect 488 239 493 277
rect 660 268 665 293
rect 698 293 828 297
rect 698 263 703 293
rect 764 239 771 271
rect 329 231 771 239
rect 824 215 828 293
rect 1031 292 1036 428
rect 1008 288 1036 292
rect 890 248 961 256
rect 823 212 841 215
rect 758 183 807 192
rect 530 150 828 154
rect 530 125 535 150
rect 489 47 554 55
rect 489 45 496 47
rect 166 36 496 45
rect 489 32 496 36
rect 495 -5 502 20
rect 154 -11 502 -5
rect 824 -82 828 150
rect 836 20 840 212
rect 951 118 961 248
rect 951 112 998 118
rect 1008 103 1012 288
rect 1204 158 1212 467
rect 1202 155 1212 158
rect 493 -88 553 -82
rect 493 -92 500 -88
rect 144 -97 500 -92
rect 493 -102 500 -97
rect 491 -141 500 -115
rect 836 -129 841 20
rect 1008 -4 1011 103
rect 1008 -7 1013 -4
rect 991 -69 998 -32
rect 888 -78 998 -69
rect 991 -79 998 -78
rect 1010 -120 1013 -7
rect 1010 -125 1016 -120
rect 821 -136 841 -129
rect 131 -145 501 -141
rect 161 -146 501 -145
rect 491 -147 500 -146
rect 821 -217 826 -136
rect 496 -224 556 -223
rect 164 -229 556 -224
rect 496 -240 503 -229
rect 1013 -234 1016 -125
rect 1202 -185 1209 155
rect 1248 53 1254 367
rect 1235 46 1258 53
rect 1202 -191 1206 -185
rect 127 -259 503 -252
rect 494 -367 557 -361
rect 494 -379 501 -367
rect 176 -390 503 -383
rect 175 -402 504 -396
rect 175 -431 182 -402
rect 1013 -471 1017 -234
rect 1235 -291 1241 46
rect 1235 -298 1243 -291
rect 1238 -299 1243 -298
rect -107 -474 1018 -471
<< metal4 >>
rect 549 552 723 559
rect 358 539 479 545
rect 787 541 794 632
rect 473 534 479 539
rect 697 536 801 541
rect 697 452 704 536
rect 601 447 704 452
rect 601 440 607 447
rect 587 436 607 440
rect 224 263 235 406
rect 587 277 592 436
rect 596 373 601 416
rect 708 373 714 374
rect 596 368 714 373
rect 487 272 592 277
rect 708 264 714 368
rect 815 277 822 407
rect 815 271 909 277
rect 708 259 718 264
rect 473 221 479 252
rect 709 228 718 259
rect 685 221 718 228
rect 473 212 694 221
rect 685 98 694 212
rect 238 90 694 98
rect 209 -47 781 -42
rect 209 -57 218 -47
rect 901 -105 909 271
rect 880 -112 910 -105
rect 315 -224 321 -204
rect 315 -230 537 -224
rect 531 -239 537 -230
rect 773 -239 779 -218
rect 531 -246 779 -239
rect 881 -274 889 -112
rect 834 -282 889 -274
rect 834 -350 843 -282
<< metal5 >>
rect 313 517 321 663
rect 702 638 778 644
rect 410 500 416 581
rect 473 529 646 533
rect 172 478 693 485
rect 513 454 639 461
rect 144 444 149 445
rect 81 441 149 444
rect 144 346 149 441
rect 702 416 708 638
rect 595 410 708 416
rect 371 407 376 408
rect 371 402 492 407
rect 826 392 837 395
rect 273 346 281 374
rect 833 351 837 392
rect 833 347 857 351
rect 144 340 282 346
rect 273 229 281 340
rect 699 327 748 333
rect 402 51 409 248
rect 448 208 455 252
rect 448 201 785 208
rect 401 37 409 51
rect 401 28 408 37
rect 401 22 409 28
rect 401 -106 408 22
rect 661 -14 667 131
rect 400 -113 408 -106
rect 400 -247 407 -113
rect 400 -286 406 -247
rect 400 -293 427 -286
rect 566 -293 573 -157
rect 758 -222 764 194
rect 776 -48 785 201
rect 849 192 856 347
rect 800 183 856 192
rect 744 -228 764 -222
rect 803 -151 809 -19
rect 400 -294 574 -293
rect 418 -301 574 -294
rect 744 -298 752 -228
rect 803 -293 812 -151
rect 418 -381 425 -301
rect 744 -356 751 -298
<< metal6 >>
rect 671 608 677 611
rect 592 603 677 608
rect 233 406 241 540
rect 313 517 314 524
rect 313 435 318 517
rect 236 395 241 406
rect 273 427 320 435
rect 273 375 282 427
rect 671 391 677 603
rect 281 369 282 375
rect 666 -126 787 -123
rect 657 -129 787 -126
rect 657 -255 666 -129
rect 793 -129 797 -123
rect 657 -256 824 -255
rect 517 -264 657 -259
rect 666 -263 819 -256
rect 517 -265 666 -264
rect 517 -274 523 -265
rect 425 -281 523 -274
rect 518 -400 523 -281
rect 668 -286 815 -285
rect 668 -290 810 -286
rect 518 -406 547 -400
rect 720 -406 812 -400
rect 518 -407 550 -406
rect 542 -459 550 -407
rect 542 -467 543 -459
<< pad >>
rect 302 655 321 662
rect 689 654 694 659
rect 722 654 727 659
rect 755 654 760 659
rect 788 654 793 659
rect 821 654 826 659
rect 208 644 216 651
rect 265 644 272 651
rect 838 646 843 651
rect 872 645 878 650
rect 772 636 778 644
rect 519 625 524 630
rect 552 625 557 630
rect 585 625 590 630
rect 618 625 623 630
rect 788 628 794 634
rect 635 617 640 622
rect 665 617 671 623
rect 382 604 387 609
rect 415 604 420 609
rect 448 604 453 609
rect 585 603 592 608
rect 465 596 470 601
rect 498 596 504 601
rect 359 591 364 596
rect 413 575 419 581
rect 573 569 581 577
rect 185 561 190 567
rect 378 561 384 567
rect 515 560 523 569
rect 401 550 407 556
rect 548 551 556 560
rect 233 540 242 547
rect 220 506 228 513
rect 172 478 178 485
rect 79 441 84 446
rect -47 420 -42 426
rect 198 410 203 415
rect 358 539 364 544
rect 249 528 255 534
rect 473 528 478 534
rect 641 529 647 534
rect 314 517 322 524
rect 277 505 284 512
rect 410 500 415 506
rect 398 462 403 467
rect 431 462 436 467
rect 464 462 469 467
rect 535 464 540 469
rect 568 464 573 469
rect 601 464 606 469
rect 634 464 639 469
rect 370 453 375 458
rect 481 454 486 459
rect 513 454 519 461
rect 636 454 642 459
rect 651 456 656 461
rect 564 440 569 445
rect 37 398 43 403
rect -116 392 -111 397
rect 225 395 236 406
rect 431 433 436 438
rect 601 436 606 441
rect -47 367 -42 373
rect 160 366 171 380
rect 531 421 536 426
rect 394 410 399 415
rect 417 408 422 413
rect 596 410 601 415
rect 371 402 378 408
rect 487 402 494 409
rect 303 390 310 397
rect 750 577 756 583
rect 684 563 692 570
rect 717 558 723 566
rect 842 494 848 501
rect 687 478 694 486
rect 1204 472 1212 479
rect 810 466 817 472
rect 867 459 873 464
rect 682 453 687 458
rect 719 454 724 459
rect 1096 451 1101 457
rect 709 444 714 449
rect 954 440 962 447
rect 871 426 876 431
rect 1180 429 1186 434
rect 1027 423 1032 428
rect 740 405 745 410
rect 774 406 779 411
rect 815 402 820 407
rect 694 394 699 399
rect 715 394 720 399
rect 744 394 749 399
rect 777 394 782 399
rect 787 394 792 399
rect 1096 398 1101 404
rect 825 392 830 397
rect 367 379 375 386
rect 671 384 677 391
rect 892 377 897 382
rect 926 379 931 384
rect 273 368 281 375
rect 330 368 337 375
rect 965 374 972 380
rect 1013 374 1019 380
rect 826 366 831 371
rect 846 366 851 371
rect 867 366 872 371
rect 896 366 901 371
rect 929 366 934 371
rect 939 366 944 371
rect 1245 361 1255 370
rect 111 333 117 340
rect 597 333 602 338
rect 834 333 842 340
rect 78 326 86 331
rect 695 327 700 332
rect 740 322 748 329
rect 425 315 430 320
rect 605 315 610 320
rect -48 306 -43 312
rect 454 301 459 306
rect 487 301 492 306
rect 520 301 525 306
rect 537 293 542 298
rect 566 293 571 298
rect 36 284 42 289
rect -117 278 -112 283
rect 487 272 493 277
rect 806 276 812 281
rect 224 263 235 271
rect 626 266 631 271
rect 660 268 665 273
rect 698 263 703 268
rect 764 265 769 271
rect -48 253 -43 259
rect 152 254 160 262
rect 601 255 606 260
rect 630 255 635 260
rect 663 255 668 260
rect 673 255 678 260
rect 714 256 723 265
rect 367 241 375 248
rect 401 241 410 248
rect 450 247 455 252
rect 473 247 478 252
rect 890 248 898 256
rect 273 230 281 237
rect 329 231 337 239
rect 812 233 818 238
rect 111 219 117 226
rect 77 213 85 218
rect -45 192 -40 198
rect 753 183 765 194
rect 800 183 809 193
rect 39 170 45 175
rect -114 164 -109 169
rect 1203 152 1208 157
rect -45 139 -40 145
rect 136 139 148 150
rect 488 130 493 135
rect 1077 131 1082 137
rect 530 125 535 130
rect 660 124 668 131
rect 332 113 337 118
rect 458 117 463 122
rect 491 117 496 122
rect 501 117 506 122
rect 566 113 574 120
rect 615 114 623 122
rect 111 105 117 112
rect 993 111 999 119
rect 1161 109 1167 114
rect 1008 103 1013 108
rect 78 98 86 103
rect 238 90 245 97
rect -42 78 -37 84
rect 381 79 386 85
rect 1077 78 1082 84
rect 337 70 343 76
rect 42 56 48 61
rect 712 58 720 66
rect 740 58 748 66
rect -111 50 -106 55
rect 554 47 562 55
rect 1235 44 1241 51
rect -42 25 -37 31
rect 125 22 137 36
rect 489 30 497 38
rect 1202 37 1210 42
rect 401 21 409 28
rect 307 10 315 17
rect 494 14 502 22
rect 1076 17 1081 23
rect 111 -9 117 -3
rect 1160 -5 1166 0
rect 657 -14 665 -7
rect 1007 -11 1012 -6
rect 83 -19 88 -14
rect 332 -21 338 -16
rect 563 -25 571 -18
rect 610 -23 617 -16
rect 803 -25 812 -18
rect -43 -40 -38 -34
rect 991 -37 1000 -28
rect 1076 -36 1081 -30
rect 776 -47 782 -41
rect 209 -57 217 -50
rect 381 -55 386 -49
rect 41 -62 47 -57
rect 337 -63 343 -58
rect -112 -68 -107 -63
rect 866 -71 872 -66
rect 1235 -70 1241 -63
rect 712 -80 720 -72
rect 741 -80 749 -72
rect 824 -82 829 -76
rect 888 -78 896 -71
rect 1201 -76 1209 -71
rect -43 -93 -38 -87
rect 552 -90 559 -83
rect 1079 -97 1084 -91
rect 401 -113 409 -106
rect 491 -108 501 -99
rect 871 -114 877 -109
rect 115 -127 121 -120
rect 307 -124 315 -117
rect 491 -124 501 -115
rect 1163 -119 1169 -114
rect 657 -126 666 -120
rect 82 -134 90 -129
rect -44 -154 -39 -148
rect 333 -155 339 -150
rect 566 -163 574 -156
rect 619 -161 626 -154
rect 40 -176 46 -171
rect -113 -182 -108 -177
rect 382 -189 387 -183
rect 338 -197 344 -192
rect -44 -207 -39 -201
rect 315 -209 321 -204
rect 153 -231 167 -219
rect 555 -229 562 -222
rect 115 -241 121 -234
rect 81 -247 89 -242
rect 400 -247 409 -240
rect 495 -244 502 -237
rect 127 -261 138 -250
rect 496 -259 503 -252
rect 787 -130 793 -123
rect 1010 -125 1015 -120
rect 1079 -150 1084 -144
rect 797 -159 805 -152
rect 1235 -184 1241 -177
rect 1202 -191 1210 -186
rect 863 -205 869 -200
rect 719 -218 724 -211
rect 743 -219 751 -211
rect 821 -216 826 -210
rect 1082 -211 1087 -205
rect 773 -224 779 -218
rect 1166 -233 1172 -228
rect 1013 -239 1018 -234
rect 869 -248 874 -243
rect -41 -268 -36 -262
rect 657 -264 666 -256
rect 819 -264 827 -256
rect 1082 -264 1087 -258
rect 419 -281 425 -273
rect 43 -290 49 -285
rect 333 -289 339 -284
rect -110 -296 -105 -291
rect -41 -321 -36 -315
rect 382 -323 387 -317
rect 338 -331 344 -326
rect 115 -355 121 -348
rect 82 -362 90 -357
rect -38 -382 -33 -376
rect 170 -386 185 -370
rect 417 -381 425 -372
rect 494 -384 501 -377
rect 46 -404 52 -399
rect 496 -400 503 -393
rect 660 -290 668 -283
rect 566 -301 574 -294
rect 617 -299 624 -292
rect 810 -293 818 -286
rect 1235 -298 1241 -292
rect 876 -339 882 -334
rect 716 -356 723 -349
rect 743 -356 751 -348
rect 834 -350 839 -344
rect 555 -367 562 -360
rect 882 -382 888 -377
rect 806 -400 812 -393
rect -107 -410 -102 -405
rect 547 -406 554 -400
rect 713 -406 720 -400
rect -38 -435 -33 -429
rect 176 -433 190 -423
rect 115 -467 121 -461
rect 543 -467 555 -459
<< labels >>
rlabel metal1 484 32 484 32 1 a0
rlabel metal1 485 15 485 15 1 b0
rlabel metal1 492 -103 492 -103 1 a1
rlabel metal1 493 -399 493 -399 1 b3
rlabel metal1 488 -121 488 -121 1 b1
rlabel metal1 418 129 418 129 5 gnd
rlabel metal1 261 79 261 79 3 p0
rlabel metal1 261 -55 261 -55 1 p1
rlabel metal1 418 -5 418 -5 5 gnd
rlabel metal1 419 -139 419 -139 5 gnd
rlabel metal1 419 -273 419 -273 5 gnd
rlabel metal1 332 237 332 237 1 cin
rlabel metal1 422 178 422 178 1 pocin
rlabel metal1 511 98 511 98 1 gnd
rlabel metal1 530 127 530 127 1 c1
rlabel metal1 424 317 424 317 1 p1g0
rlabel metal1 451 292 451 292 1 p1
rlabel metal1 475 292 475 292 1 p0
rlabel metal1 489 285 489 285 1 cin
rlabel metal1 211 405 211 405 1 gnd
rlabel metal1 489 388 489 388 1 gnd
rlabel metal1 533 443 533 443 1 p2
rlabel metal1 565 446 565 446 1 p1
rlabel metal1 589 447 589 447 1 p0
rlabel metal1 602 442 602 442 1 cin
rlabel metal1 680 458 680 458 1 p2p1p0c0
rlabel metal1 691 407 691 407 1 g2
rlabel pad 742 408 742 408 1 p2p1p0c0
rlabel metal1 202 444 202 444 3 p2
rlabel metal1 368 454 368 454 1 p2g1
rlabel metal1 396 449 396 449 1 p2
rlabel metal1 418 449 418 449 1 p1
rlabel metal1 434 441 434 441 1 g0
rlabel metal1 511 457 511 457 1 p2p1g0
rlabel metal1 775 409 775 409 1 p2g1
rlabel metal1 199 543 199 543 1 gnd
rlabel metal1 473 530 473 530 1 gnd
rlabel metal1 643 551 643 551 1 gnd
rlabel metal1 192 583 192 583 1 p3
rlabel metal1 264 652 264 652 1 g2
rlabel metal1 359 593 359 593 1 p3g2
rlabel metal1 379 591 379 591 1 p3
rlabel metal1 402 591 402 591 1 p2
rlabel metal1 418 585 418 585 1 g1
rlabel metal1 494 597 494 597 1 p3p2g1
rlabel metal1 516 599 516 599 1 p3
rlabel metal1 550 603 550 603 1 p2
rlabel metal1 586 604 586 604 1 g0
rlabel metal1 666 619 666 619 1 p3p2p1g0
rlabel metal1 686 633 686 633 1 p3
rlabel metal1 720 624 720 624 1 p2
rlabel metal1 753 631 753 631 1 p1
rlabel metal1 775 638 775 638 1 p0
rlabel metal1 790 636 790 636 1 cin
rlabel metal1 867 648 867 648 1 p3p2p1p0c0
rlabel metal1 824 398 824 398 1 g3
rlabel metal1 843 395 843 395 1 p3g2
rlabel metal1 864 395 864 395 1 p3p2g1
rlabel metal1 928 379 928 379 1 p3p2p1p0c0
rlabel metal1 726 260 726 260 1 p0
rlabel pad 766 268 766 268 1 cin
rlabel pad 894 380 894 380 1 p3p2p1g0
rlabel metal1 570 295 570 295 1 p1p0c0
rlabel pad 489 131 489 131 1 g0
rlabel metal1 698 265 698 265 1 c2
rlabel metal1 598 272 598 272 1 g1
rlabel pad 628 267 628 267 1 p1g0
rlabel metal1 661 268 661 268 1 p1p0c0
rlabel metal1 573 612 573 612 1 p1
rlabel metal1 712 409 712 409 1 p2p1g0
rlabel metal1 316 -322 316 -322 1 p3
rlabel metal1 319 -189 319 -189 1 p2
rlabel metal1 815 404 815 404 7 c3
rlabel metal1 483 -257 483 -257 1 b2
rlabel metal1 619 14 619 14 1 gnd
rlabel metal1 757 62 757 62 1 g0
rlabel metal1 554 -126 554 -126 1 gnd
rlabel metal1 557 -264 557 -264 1 gnd
rlabel metal1 557 -402 557 -402 1 gnd
rlabel metal1 836 -343 836 -343 1 c3
rlabel pad 836 -348 836 -348 1 c3
rlabel metal1 791 -356 791 -356 1 p3
rlabel metal1 801 -394 801 -394 1 gnd
rlabel pad 823 -213 823 -213 1 c2
rlabel metal1 777 -221 777 -221 1 p2
rlabel metal1 788 -260 788 -260 1 gnd
rlabel metal1 761 -212 761 -212 1 g2
rlabel metal1 783 -87 783 -87 1 p1
rlabel pad 825 -79 825 -79 1 c1
rlabel metal1 269 514 269 514 1 g1
rlabel metal1 751 -76 751 -76 1 g1
rlabel metal1 762 -353 762 -353 1 g3
rlabel metal1 -76 364 -76 364 7 gnd
rlabel metal1 -6 364 -6 364 7 gnd
rlabel metal1 -118 394 -118 394 3 clk
rlabel metal1 56 364 56 364 7 gnd
rlabel metal1 98 335 98 335 1 gnd
rlabel metal1 97 221 97 221 1 gnd
rlabel metal1 55 250 55 250 7 gnd
rlabel metal1 -119 280 -119 280 3 clk
rlabel metal1 -7 250 -7 250 7 gnd
rlabel metal1 -77 250 -77 250 7 gnd
rlabel metal1 100 107 100 107 1 gnd
rlabel metal1 58 136 58 136 7 gnd
rlabel metal1 -116 166 -116 166 3 clk
rlabel metal1 -4 136 -4 136 7 gnd
rlabel metal1 -74 136 -74 136 7 gnd
rlabel metal1 -71 22 -71 22 7 gnd
rlabel metal1 -1 22 -1 22 7 gnd
rlabel metal1 -113 52 -113 52 3 clk
rlabel metal1 61 22 61 22 7 gnd
rlabel metal1 103 -7 103 -7 1 gnd
rlabel metal1 -72 -96 -72 -96 7 gnd
rlabel metal1 -2 -96 -2 -96 7 gnd
rlabel metal1 -114 -66 -114 -66 3 clk
rlabel metal1 60 -96 60 -96 7 gnd
rlabel metal1 102 -125 102 -125 1 gnd
rlabel metal1 101 -239 101 -239 1 gnd
rlabel metal1 59 -210 59 -210 7 gnd
rlabel metal1 -115 -180 -115 -180 3 clk
rlabel metal1 -3 -210 -3 -210 7 gnd
rlabel metal1 -73 -210 -73 -210 7 gnd
rlabel metal1 104 -353 104 -353 1 gnd
rlabel metal1 62 -324 62 -324 7 gnd
rlabel metal1 -112 -294 -112 -294 3 clk
rlabel metal1 0 -324 0 -324 7 gnd
rlabel metal1 -70 -324 -70 -324 7 gnd
rlabel metal1 -67 -438 -67 -438 7 gnd
rlabel metal1 3 -438 3 -438 7 gnd
rlabel metal1 -109 -408 -109 -408 3 clk
rlabel metal1 65 -438 65 -438 7 gnd
rlabel metal1 107 -467 107 -467 1 gnd
rlabel metal1 -127 397 -127 397 3 a0_in
rlabel metal1 -128 297 -128 297 3 b0_in
rlabel metal1 -125 181 -125 181 3 a1_in
rlabel metal1 -122 54 -122 54 1 b1_in
rlabel metal1 -124 -173 -124 -173 3 b2_in
rlabel metal1 -121 -297 -121 -297 1 a3_in
rlabel metal1 -118 -403 -118 -403 1 b3_in
rlabel metal1 125 -431 125 -431 1 b3
rlabel metal1 124 -203 124 -203 1 b2
rlabel metal1 118 29 118 29 1 b1
rlabel metal1 111 370 111 370 1 a0
rlabel metal1 1067 395 1067 395 7 gnd
rlabel metal1 1137 395 1137 395 7 gnd
rlabel metal1 1025 425 1025 425 3 clk
rlabel metal1 1199 395 1199 395 7 gnd
rlabel metal1 1241 366 1241 366 1 gnd
rlabel metal1 1048 75 1048 75 7 gnd
rlabel metal1 1118 75 1118 75 7 gnd
rlabel metal1 1006 105 1006 105 3 clk
rlabel metal1 1180 75 1180 75 7 gnd
rlabel metal1 1222 46 1222 46 1 gnd
rlabel metal1 1221 -68 1221 -68 1 gnd
rlabel metal1 1179 -39 1179 -39 7 gnd
rlabel metal1 1005 -9 1005 -9 3 clk
rlabel metal1 1117 -39 1117 -39 7 gnd
rlabel metal1 1047 -39 1047 -39 7 gnd
rlabel metal1 1224 -182 1224 -182 1 gnd
rlabel metal1 1182 -153 1182 -153 7 gnd
rlabel metal1 1008 -123 1008 -123 3 clk
rlabel metal1 1120 -153 1120 -153 7 gnd
rlabel metal1 1050 -153 1050 -153 7 gnd
rlabel metal1 1053 -267 1053 -267 7 gnd
rlabel metal1 1123 -267 1123 -267 7 gnd
rlabel metal1 1011 -237 1011 -237 3 clk
rlabel metal1 1185 -267 1185 -267 7 gnd
rlabel metal1 1227 -296 1227 -296 1 gnd
rlabel metal1 950 347 950 347 1 gnd
rlabel metal1 732 221 732 221 1 gnd
rlabel metal1 792 -126 792 -126 1 gnd
rlabel metal1 546 227 546 227 1 gnd
rlabel metal1 419 267 419 267 5 gnd
rlabel metal1 684 236 684 236 1 gnd
rlabel metal1 798 375 798 375 1 gnd
rlabel metal1 660 390 660 390 1 gnd
rlabel metal1 847 580 847 580 1 gnd
rlabel metal1 962 376 962 376 1 c4_in
rlabel metal1 493 -243 493 -243 1 a2
rlabel metal1 894 269 894 269 1 s0_in
rlabel metal1 1253 402 1253 402 7 c4
rlabel metal1 1233 -32 1233 -32 1 s1
rlabel metal1 1232 -146 1232 -146 1 s2
rlabel metal1 1243 -259 1243 -259 1 s3
rlabel pad 892 -75 892 -75 1 s1_in
rlabel metal1 902 -343 902 -343 1 s3_in
rlabel metal1 890 -210 890 -210 1 s2_in
rlabel metal1 1245 474 1245 474 5 vdd
rlabel metal1 803 470 803 470 5 vdd
rlabel metal1 1226 154 1226 154 5 vdd
rlabel metal1 1228 -74 1228 -74 5 vdd
rlabel metal1 1225 40 1225 40 5 vdd
rlabel metal1 1231 -188 1231 -188 5 vdd
rlabel metal1 955 442 955 442 5 vdd
rlabel metal1 689 331 689 331 5 vdd
rlabel metal1 507 363 507 363 5 vdd
rlabel metal1 378 381 378 381 5 vdd
rlabel metal1 411 381 411 381 5 vdd
rlabel metal1 204 646 204 646 5 vdd
rlabel metal1 346 657 346 657 5 vdd
rlabel metal1 435 666 435 666 5 vdd
rlabel metal1 605 687 605 687 5 vdd
rlabel metal1 808 716 808 716 5 vdd
rlabel metal1 216 508 216 508 5 vdd
rlabel metal1 358 519 358 519 5 vdd
rlabel metal1 451 524 451 524 5 vdd
rlabel metal1 621 526 621 526 5 vdd
rlabel metal1 378 243 378 243 5 vdd
rlabel metal1 411 243 411 243 5 vdd
rlabel metal1 414 -242 414 -242 1 vdd
rlabel metal1 793 -157 793 -157 5 vdd
rlabel metal1 800 -23 800 -23 5 vdd
rlabel metal1 806 -291 806 -291 5 vdd
rlabel metal1 704 -288 704 -288 5 vdd
rlabel metal1 671 -288 671 -288 5 vdd
rlabel metal1 562 -299 562 -299 5 vdd
rlabel metal1 414 -376 414 -376 1 vdd
rlabel metal1 562 -161 562 -161 5 vdd
rlabel metal1 304 -119 304 -119 1 vdd
rlabel metal1 413 -108 413 -108 1 vdd
rlabel metal1 304 15 304 15 1 vdd
rlabel metal1 413 26 413 26 1 vdd
rlabel metal1 517 193 517 193 5 vdd
rlabel metal1 704 126 704 126 5 vdd
rlabel metal1 671 126 671 126 5 vdd
rlabel metal1 559 -23 559 -23 5 vdd
rlabel metal1 668 -12 668 -12 5 vdd
rlabel metal1 701 -12 701 -12 5 vdd
rlabel metal1 562 115 562 115 5 vdd
rlabel metal1 269 232 269 232 5 vdd
rlabel metal1 104 215 104 215 5 vdd
rlabel metal1 101 329 101 329 5 vdd
rlabel metal1 107 101 107 101 5 vdd
rlabel metal1 111 -359 111 -359 5 vdd
rlabel metal1 108 -245 108 -245 5 vdd
rlabel metal1 105 -131 105 -131 5 vdd
rlabel metal1 106 -17 106 -17 5 vdd
rlabel metal1 102 443 102 443 5 vdd
rlabel metal1 269 370 269 370 5 vdd
rlabel metal1 736 324 736 324 5 vdd
rlabel metal1 878 335 878 335 5 vdd
rlabel metal1 845 335 845 335 5 vdd
rlabel metal1 -123 -54 -123 -54 1 a2_in
rlabel metal1 484 -383 484 -383 1 a3
rlabel metal1 123 -317 123 -317 1 a3
rlabel metal1 1235 82 1235 82 1 s0
rlabel metal1 121 -89 121 -89 1 a2
rlabel metal1 125 144 125 144 1 a1
rlabel metal1 122 256 122 256 1 b0
<< end >>
