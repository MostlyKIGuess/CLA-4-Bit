* SPICE3 file created from testing.ext - technology: scmos

.option scale=1u

M1000 g2 a_582_n251# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 a_445_147# g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 p2g1 a_327_429# vdd w_347_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1003 a_594_575# p1 a_594_556# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_440_412# p1 a_440_393# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1005 p1p0c0 a_453_311# vdd w_544_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 a3 b3 p3 w_329_n384# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 s2 p2 c2 w_835_n8# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 a_518_635# p3 vdd w_505_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1009 a_731_457# p2p1p0c0 a_731_417# w_725_444# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 b2 a2 p2 w_368_n246# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1011 p3p2g1 a_381_614# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 p2p1p0c0 a_534_474# vdd w_658_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1013 a_610_395# p1 a_610_377# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1014 b2 a_325_n180# p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1015 a_815_n46# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1016 a_518_635# g0 a_594_575# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1017 vdd a0 a_324_88# w_400_28# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1018 vdd a_302_20# a_269_20# w_291_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_325_n180# b2 p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1020 g0 a_691_36# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1021 a_825_350# p3p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1022 a_304_190# a_271_142# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1023 a_847_245# a_771_282# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1024 a_884_498# p3g2 a_883_464# w_878_485# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1025 g3 a_691_n378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1026 a_731_492# p2p1g0 a_731_457# w_725_479# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1027 s1 a_798_100# c1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1028 a_615_n341# a3 b3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1029 a_798_100# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 s1 c1 p1 w_857_146# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 a_315_567# a_239_604# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 a_582_n251# a2 vdd w_569_n219# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1033 p3g2 a_315_567# vdd w_335_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1034 vdd g3 a_884_498# w_879_518# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 a_825_350# p3p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 pocin a_380_153# vdd w_400_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1037 vdd a_269_20# p0 w_258_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1038 a_218_418# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1039 a_380_153# a_304_190# vdd w_367_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 b1 a1 a_302_n114# w_367_n112# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1041 a_691_36# a_615_73# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 a_825_350# p3p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1043 a_271_280# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 p3p2p1g0 a_518_635# vdd w_642_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 g2 a_582_n251# b2 w_602_n213# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 a_239_604# a_206_556# g2 w_226_594# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1047 a_304_190# a_271_142# cin w_291_180# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1048 a_612_n65# a_579_n113# b1 w_599_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 a_582_25# a0 vdd w_569_57# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 p2p1g0 a_397_472# vdd w_488_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1051 c3 a_693_378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1052 a_440_393# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_612_n65# a_579_n113# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1054 a_688_664# p0 vdd w_774_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1055 a_445_147# pocin gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1056 p2g1 a_327_429# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1057 a_600_239# p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1058 a_327_429# a_251_466# vdd w_314_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1059 s2 a_815_n46# c2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 a_688_664# cin vdd w_807_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_693_378# p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1062 a_251_466# p2 g1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1063 a_325_n314# b3 p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1064 a_688_n102# a_612_n65# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 a_738_234# p0 vdd w_725_266# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1066 p3p2g1 a_381_614# vdd w_472_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1067 a_206_556# p3 vdd w_193_588# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_424_535# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_610_377# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 s0 a_847_245# vdd w_867_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1071 a_582_n389# a3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_691_n378# a_615_n341# vdd w_678_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1073 s3 a_831_n180# c3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 vdd a2 a_325_n180# w_401_n240# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 g2 a2 b2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 g1 a_688_n102# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1077 c4 a_825_350# vdd w_942_382# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1078 a_424_554# p2 a_424_535# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1079 a_453_311# p0 vdd w_473_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1080 a_831_n180# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1081 a_315_567# a_239_604# vdd w_302_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 p3p2p1p0c0 a_688_664# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1083 a_771_282# p0 cin w_758_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1084 a_612_n65# a1 b1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1085 a_271_142# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1086 a_534_474# cin vdd w_620_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1087 a_534_474# p0 vdd w_587_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1088 a_453_311# cin vdd w_506_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_271_280# p1 vdd w_258_312# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 a_693_378# p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1091 a_381_614# g1 a_424_554# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1092 a_883_429# p3p2p1g0 a_883_389# w_877_416# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 c1 a_445_147# vdd w_504_133# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1094 a_304_328# a_271_280# g0 w_291_318# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 a_825_350# p3g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_688_664# p1 vdd w_741_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1097 a_797_604# p0 a_797_585# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 vdd a_269_n114# p1 w_258_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1099 p1g0 a_380_291# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1100 a_324_n46# b1 a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1101 a_327_429# a_251_466# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1102 a1 b1 a_302_n114# w_328_n116# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_693_378# p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1104 a_380_291# a_304_328# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1105 c2 a_600_239# vdd w_676_271# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 b3 a3 p3 w_368_n380# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1107 a_688_n102# a_612_n65# vdd w_675_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 b1 a_324_n46# a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1109 a_815_n46# p2 vdd w_802_n14# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1110 b0 a_324_88# a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 vdd a3 a_325_n314# w_401_n374# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1112 a_615_73# a_582_25# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1113 p1p0c0 a_453_311# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1114 a_324_88# b0 a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1115 a_688_664# cin a_797_604# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1116 vdd g2 a_731_492# w_726_513# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1117 a_883_464# p3p2g1 a_883_429# w_877_451# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1118 a_693_378# g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 g1 a_688_n102# vdd w_708_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1120 s1 c1 a_798_100# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1121 s3 p3 c3 w_851_n142# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1122 a_304_328# p1 g0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1123 a_771_282# a_738_234# cin Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1124 a_518_635# p1 vdd w_571_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1125 a_397_472# g0 vdd w_450_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1126 a_579_n113# a1 vdd w_566_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1127 a_797_547# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1128 a_496_251# p0 a_496_232# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1129 s2 c2 p2 w_874_0# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 a_518_635# g0 vdd w_604_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1131 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 p2p1p0c0 a_534_474# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 g0 a_691_36# vdd w_711_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1134 a_847_245# a_771_282# vdd w_834_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1135 a_579_n113# a1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1136 a_239_604# a_206_556# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1137 a_797_566# p2 a_797_547# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1138 a_453_311# cin a_496_251# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_453_311# p1 vdd w_440_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 gnd a3 a_325_n314# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1141 a_798_100# p1 vdd w_785_132# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_534_474# p1 vdd w_554_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_304_328# a_271_280# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1144 a_445_147# g0 a_445_140# w_439_134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1145 a_797_585# p1 a_797_566# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 s3 c3 a_831_n180# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1147 gnd a_302_n114# a_269_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1148 a_691_36# a_615_73# vdd w_678_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1149 s3 c3 p3 w_890_n134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1150 gnd a_269_n114# p1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1151 a_381_614# g1 vdd w_434_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1152 s2 c2 a_815_n46# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1153 pocin a_380_153# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1154 s1 p1 c1 w_818_138# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 a_380_153# a_304_190# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1156 a_688_664# p3 vdd w_675_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1157 g3 a_691_n378# vdd w_711_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1158 p1g0 a_380_291# vdd w_400_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1159 c2 a_600_239# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1160 a0 b0 a_302_20# w_328_18# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 a_615_73# a0 b0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_380_291# a_304_328# vdd w_367_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1163 a_582_25# a0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_688_664# p2 vdd w_708_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1165 p2p1g0 a_397_472# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1166 gnd a2 a_325_n180# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1167 vdd pocin a_445_140# w_439_167# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 c3 a_693_378# vdd w_790_410# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1169 a_304_190# p0 cin Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1170 a_251_466# a_218_418# g1 w_238_456# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1171 vdd a1 a_324_n46# w_400_n106# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1172 a_397_472# g0 a_440_412# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 a_691_n378# a_615_n341# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1174 a_615_n341# a_582_n389# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1175 a_397_472# p2 vdd w_384_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1176 vdd a_302_n114# a_269_n114# w_291_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1177 a_617_318# p1g0 a_617_278# w_611_305# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1178 a_771_282# cin p0 w_797_280# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_738_234# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1180 a_518_635# p2 vdd w_538_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1181 b0 a0 a_302_20# w_367_22# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1182 a_496_232# p1 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 a_397_472# p1 vdd w_417_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1184 a_206_556# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1185 a_610_414# p0 a_610_395# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 p3p2p1p0c0 a_688_664# vdd w_845_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1187 a_271_142# p0 vdd w_258_174# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1188 a_582_n251# a2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1189 a_534_474# p2 vdd w_521_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 s0 a_847_245# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1191 vdd g1 a_617_318# w_611_340# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1192 c4 a_825_350# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1193 gnd a1 a_324_n46# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1194 gnd a0 a_324_88# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1195 gnd a_302_20# a_269_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1196 a_381_614# p2 vdd w_401_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 a_534_474# cin a_610_414# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a2 b2 p2 w_329_n250# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1199 a_251_466# a_218_418# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1200 a_771_282# cin a_738_234# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1201 a_381_614# p3 vdd w_368_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 p3g2 a_315_567# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1203 a_594_537# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_600_239# g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1205 a_615_73# a_582_25# b0 w_602_63# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1206 a_582_n389# a3 vdd w_569_n357# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 a_239_604# p3 g2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1208 b3 a_325_n314# p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1209 a_218_418# p2 vdd w_205_450# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1210 a_825_350# g3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1211 a_600_239# p1p0c0 a_617_278# w_611_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1212 c1 a_445_147# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1213 p3p2p1g0 a_518_635# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 a_693_378# p2g1 a_731_417# w_725_411# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1215 a_831_n180# p3 vdd w_818_n148# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1216 a_600_239# p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1217 a_594_556# p2 a_594_537# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1218 gnd a_269_20# p0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1219 a_615_n341# a_582_n389# b3 w_602_n351# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 w_818_138# s1 2.162f
C1 w_675_654# a_688_664# 2.45f
C2 w_400_323# a_380_291# 1.014f
C3 a_534_474# p1 0.19f
C4 w_725_266# vdd 1.128f
C5 w_488_462# vdd 1.128f
C6 a_397_472# p1 0.19f
C7 w_329_n384# p3 1.128f
C8 w_802_n14# a_815_n46# 1.88f
C9 w_571_625# a_518_635# 3.59f
C10 w_401_n240# a2 1.014f
C11 w_314_461# a_251_466# 1.014f
C12 g1 gnd 15.03f
C13 w_472_604# a_381_614# 1.014f
C14 w_400_323# g0 1.33f
C15 w_890_n134# s3 1.128f
C16 w_521_464# p2 1.014f
C17 w_818_138# c1 1.88f
C18 g0 a_380_291# 1.01f
C19 w_384_462# vdd 1.128f
C20 w_790_410# c3 1.88f
C21 g1 vdd 2.472f
C22 a_381_614# p2 0.19f
C23 w_368_604# a_381_614# 2.45f
C24 w_878_485# a_883_464# 1.41f
C25 w_711_68# vdd 1.128f
C26 w_226_594# a_206_556# 1.014f
C27 w_473_301# p0 1.014f
C28 a_534_474# cin 0.19f
C29 w_890_n134# c3 1.17f
C30 w_506_301# vdd 1.128f
C31 w_878_485# p3g2 1.482f
C32 w_818_138# p1 1.17f
C33 a_304_328# g0 1.35f
C34 a_518_635# p2 0.19f
C35 a_534_474# p0 0.19f
C36 w_890_n134# p3 1.128f
C37 w_802_n14# p2 1.014f
C38 w_439_134# a_445_140# 2.444f
C39 w_678_n346# vdd 1.128f
C40 b0 a_302_20# 4.68f
C41 w_571_625# p1 1.014f
C42 a_688_664# p2 0.19f
C43 w_569_57# vdd 1.128f
C44 w_439_134# a_445_147# 1.88f
C45 w_797_280# a_771_282# 1.128f
C46 w_604_625# g0 1.014f
C47 w_400_323# vdd 1.128f
C48 w_226_594# a_239_604# 2.82f
C49 w_676_271# a_600_239# 1.014f
C50 w_774_654# p0 1.014f
C51 w_807_654# vdd 1.128f
C52 w_678_n346# a_691_n378# 1.88f
C53 w_335_599# p3g2 1.88f
C54 b0 a_324_88# 2.925f
C55 w_504_133# g0 1.33f
C56 w_401_n374# vdd 1.128f
C57 w_602_63# a_582_25# 1.014f
C58 w_258_312# vdd 1.128f
C59 w_708_n70# a_688_n102# 1.014f
C60 g0 vdd 4.29f
C61 a0 b0 4.458f
C62 w_708_654# vdd 1.128f
C63 w_877_416# a_883_389# 1.128f
C64 w_488_462# p2p1g0 1.88f
C65 a_304_328# vdd 1.89f
C66 w_401_n374# a_325_n314# 1.88f
C67 w_877_416# p3p2p1g0 1.482f
C68 w_566_n81# a_579_n113# 1.88f
C69 w_678_n346# a_615_n341# 1.014f
C70 w_587_464# a_534_474# 3.59f
C71 w_878_485# a_884_498# 1.598f
C72 w_193_588# p3 1.014f
C73 w_401_n374# b3 1.71f
C74 w_726_513# a_731_492# 1.41f
C75 w_604_625# vdd 1.128f
C76 w_611_340# a_617_318# 1.41f
C77 a_615_73# b0 1.91f
C78 w_367_185# a_380_153# 1.88f
C79 w_401_n374# a3 1.014f
C80 w_726_513# g2 1.482f
C81 w_367_22# a_302_20# 2.162f
C82 w_611_340# g1 1.482f
C83 w_504_133# vdd 1.128f
C84 w_602_63# b0 1.128f
C85 a_825_350# gnd 3.232f
C86 w_505_625# vdd 1.128f
C87 w_488_462# a_397_472# 1.014f
C88 w_725_411# p2g1 2.202f
C89 w_328_n116# a_302_n114# 1.128f
C90 c1 s1 4.68f
C91 w_400_185# vdd 1.128f
C92 a_218_418# g1 1.212f
C93 w_367_22# b0 1.88f
C94 w_193_588# g2 1.064f
C95 w_538_625# p2 1.014f
C96 w_205_450# g1 1.596f
C97 w_258_n117# p1 1.88f
C98 w_258_17# a_269_20# 1.014f
C99 g1 p3 83.43f
C100 c1 a_798_100# 1.845f
C101 w_473_301# a_453_311# 3.59f
C102 w_367_22# a0 1.17f
C103 w_401_604# vdd 1.128f
C104 b3 gnd 1.73f
C105 w_602_n213# a_582_n251# 1.014f
C106 w_384_462# a_397_472# 2.45f
C107 w_602_63# a_615_73# 2.82f
C108 w_620_464# cin 1.014f
C109 w_417_462# p1 1.014f
C110 w_675_n70# vdd 1.128f
C111 w_877_416# a_883_429# 1.41f
C112 w_238_456# a_218_418# 1.014f
C113 w_845_654# a_688_664# 1.014f
C114 w_450_462# g0 1.014f
C115 w_725_411# a_731_417# 2.444f
C116 w_258_174# vdd 1.128f
C117 w_367_185# a_304_190# 1.014f
C118 w_566_n81# a1 1.014f
C119 a_518_635# p1 0.19f
C120 w_658_464# vdd 1.128f
C121 w_867_277# s0 1.88f
C122 w_602_n213# b2 1.128f
C123 b3 vdd 0.72f
C124 w_758_272# cin 1.88f
C125 w_302_599# vdd 1.128f
C126 a_688_664# p1 0.19f
C127 a3 vdd 2.52f
C128 w_400_n106# vdd 1.128f
C129 w_328_n116# b1 1.17f
C130 w_741_654# a_688_664# 3.59f
C131 w_758_272# p0 1.17f
C132 w_874_0# s2 1.128f
C133 g2 g1 2.97f
C134 a_615_n341# vdd 1.08f
C135 w_328_n116# a1 1.128f
C136 w_554_464# vdd 1.128f
C137 a_693_378# gnd 2.424f
C138 w_368_n246# b2 1.88f
C139 w_642_625# a_518_635# 1.014f
C140 w_440_301# p1 1.014f
C141 b2 gnd 1.91f
C142 b3 a_325_n314# 2.925f
C143 w_725_411# a_693_378# 1.88f
C144 w_291_n117# vdd 1.128f
C145 a_251_466# g1 1.212f
C146 w_367_323# a_380_291# 1.88f
C147 w_676_271# vdd 1.128f
C148 w_942_382# c4 1.88f
C149 w_785_132# a_798_100# 1.88f
C150 w_450_462# vdd 1.128f
C151 a3 b3 3.738f
C152 w_658_464# p2p1p0c0 1.88f
C153 w_538_625# a_518_635# 3.59f
C154 w_368_n246# a2 1.17f
C155 a_688_664# cin 0.19f
C156 a_397_472# g0 0.19f
C157 w_238_456# a_251_466# 2.82f
C158 w_434_604# a_381_614# 3.59f
C159 w_367_323# g0 1.33f
C160 w_741_654# p1 1.014f
C161 a_615_n341# b3 1.91f
C162 w_851_n142# s3 2.162f
C163 g1 a1 16.199999f
C164 w_725_479# a_731_457# 1.41f
C165 a_688_664# p0 0.19f
C166 w_611_340# vdd 1.88f
C167 w_874_0# c2 1.17f
C168 w_367_323# a_304_328# 1.014f
C169 w_347_461# vdd 1.128f
C170 w_335_599# a_315_567# 1.014f
C171 w_725_479# p2p1g0 1.482f
C172 w_874_0# p2 1.128f
C173 w_867_277# a_847_245# 1.014f
C174 a2 vdd 2.52f
C175 w_678_68# vdd 1.128f
C176 w_347_461# p2g1 1.88f
C177 w_193_588# a_206_556# 1.88f
C178 w_384_462# p2 1.014f
C179 w_611_272# p1p0c0 2.202f
C180 w_851_n142# c3 1.88f
C181 w_473_301# vdd 1.128f
C182 w_505_625# p3 1.014f
C183 g1 p2 3.825f
C184 w_602_n213# g2 2.82f
C185 w_785_132# p1 1.014f
C186 w_205_450# vdd 1.128f
C187 w_611_272# a_617_278# 2.444f
C188 w_851_n142# p3 1.17f
C189 w_439_167# a_445_140# 1.128f
C190 w_400_28# vdd 1.128f
C191 w_544_301# p1p0c0 1.88f
C192 w_758_272# a_771_282# 2.162f
C193 w_602_n351# a_582_n389# 1.014f
C194 w_367_323# vdd 1.128f
C195 w_611_272# a_600_239# 1.88f
C196 w_711_68# a_691_36# 1.014f
C197 w_774_654# vdd 1.128f
C198 g2 gnd 19.485f
C199 w_439_134# g0 2.943f
C200 b2 a_325_n180# 2.925f
C201 w_439_167# pocin 1.482f
C202 w_258_17# p0 1.88f
C203 w_291_17# vdd 1.128f
C204 w_569_57# a_582_25# 1.88f
C205 p3 b3 4.68f
C206 w_658_464# a_534_474# 1.014f
C207 w_942_382# vdd 1.128f
C208 g2 vdd 2.068f
C209 w_602_n351# b3 1.128f
C210 w_942_382# a_825_350# 1.014f
C211 w_725_479# a_731_492# 1.598f
C212 w_675_n70# a_688_n102# 1.88f
C213 w_675_654# vdd 1.128f
C214 w_569_n219# vdd 1.128f
C215 a_381_614# g1 0.19f
C216 b1 gnd 2.314f
C217 w_708_654# p2 1.014f
C218 a_251_466# vdd 1.89f
C219 w_602_n351# a_615_n341# 2.82f
C220 w_554_464# a_534_474# 3.59f
C221 w_291_180# a_271_142# 1.014f
C222 w_368_n380# b3 1.88f
C223 a2 b2 3.468f
C224 w_571_625# vdd 1.128f
C225 w_368_n380# a3 1.17f
C226 b1 vdd 0.9f
C227 w_328_18# a_302_20# 1.128f
C228 a_738_234# cin 1.845f
C229 a1 vdd 2.52f
C230 c3 s3 4.68f
C231 w_544_301# a_453_311# 1.014f
C232 w_368_n246# p2 2.162f
C233 w_569_57# a0 1.014f
C234 w_472_604# vdd 1.128f
C235 w_291_180# cin 1.128f
C236 a_612_n65# vdd 1.35f
C237 w_450_462# a_397_472# 3.59f
C238 c3 a_831_n180# 1.845f
C239 w_400_n106# a_324_n46# 1.88f
C240 g2 a_615_n341# 1.485f
C241 w_818_n148# vdd 1.128f
C242 w_291_n117# a_302_n114# 1.014f
C243 w_879_518# g3 1.482f
C244 w_367_185# vdd 1.128f
C245 w_328_18# b0 1.17f
C246 w_291_n117# a_269_n114# 1.88f
C247 w_879_518# vdd 1.88f
C248 w_440_301# a_453_311# 2.45f
C249 w_328_18# a0 1.128f
C250 w_368_604# vdd 1.128f
C251 w_569_n219# a_582_n251# 1.88f
C252 w_675_n70# a_612_n65# 1.014f
C253 w_877_451# a_883_429# 1.41f
C254 w_400_n106# b1 1.71f
C255 w_205_450# a_218_418# 1.88f
C256 w_807_654# a_688_664# 3.59f
C257 g2 b2 1.91f
C258 w_725_444# a_731_417# 1.128f
C259 w_867_277# vdd 1.128f
C260 w_347_461# a_327_429# 1.014f
C261 w_291_180# a_304_190# 2.82f
C262 w_401_604# p2 1.014f
C263 w_587_464# p0 1.014f
C264 w_877_451# p3p2g1 1.482f
C265 w_400_n106# a1 1.014f
C266 w_620_464# vdd 1.128f
C267 w_725_444# p2p1p0c0 1.482f
C268 a_518_635# g0 0.19f
C269 w_291_318# a_271_280# 1.014f
C270 w_845_654# p3p2p1p0c0 1.88f
C271 w_708_654# a_688_664# 3.59f
C272 w_857_146# s1 1.128f
C273 w_725_266# p0 1.014f
C274 w_835_n8# s2 2.162f
C275 b0 gnd 1.91f
C276 a_771_282# cin 4.68f
C277 w_521_464# vdd 1.128f
C278 w_329_n250# b2 1.17f
C279 w_368_n380# p3 2.162f
C280 w_472_604# p3p2g1 1.88f
C281 w_604_625# a_518_635# 3.59f
C282 g0 c1 1.01f
C283 w_569_n219# a2 1.014f
C284 w_725_266# a_738_234# 1.88f
C285 w_258_n117# vdd 1.128f
C286 w_877_451# a_883_464# 1.598f
C287 b0 vdd 0.9f
C288 g2 p3 1.575f
C289 w_725_444# a_731_457# 1.41f
C290 w_857_146# c1 1.17f
C291 w_675_654# p3 1.014f
C292 a0 vdd 2.52f
C293 w_417_462# vdd 1.128f
C294 w_676_271# c2 1.88f
C295 a_453_311# cin 0.19f
C296 g0 a_445_147# 0.72f
C297 a_239_604# vdd 1.89f
C298 w_505_625# a_518_635# 2.45f
C299 w_506_301# cin 1.014f
C300 w_258_312# p1 1.014f
C301 w_877_383# p3p2p1p0c0 2.202f
C302 w_329_n250# a2 1.128f
C303 w_401_604# a_381_614# 3.59f
C304 a_453_311# p0 0.19f
C305 w_291_318# g0 1.128f
C306 w_802_n14# vdd 1.128f
C307 w_544_301# vdd 1.128f
C308 p2 b2 4.68f
C309 w_835_n8# c2 1.88f
C310 w_504_133# c1 1.88f
C311 w_291_318# a_304_328# 2.82f
C312 w_711_n346# g3 1.88f
C313 w_818_n148# a_831_n180# 1.88f
C314 w_434_604# g1 1.014f
C315 w_857_146# p1 1.128f
C316 w_314_461# vdd 1.128f
C317 w_302_599# a_315_567# 1.88f
C318 w_835_n8# p2 1.17f
C319 a_615_73# vdd 1.35f
C320 w_708_n70# g1 1.88f
C321 w_834_277# a_847_245# 1.88f
C322 w_711_n346# vdd 1.128f
C323 w_807_654# cin 1.014f
C324 a_445_147# gnd 0.808f
C325 w_504_133# a_445_147# 1.014f
C326 w_834_277# a_771_282# 1.014f
C327 w_440_301# vdd 1.128f
C328 w_302_599# a_239_604# 1.014f
C329 w_845_654# vdd 1.128f
C330 w_611_305# a_617_278# 1.128f
C331 w_711_n346# a_691_n378# 1.014f
C332 w_818_n148# p3 1.014f
C333 w_569_n357# vdd 1.128f
C334 b1 a_302_n114# 4.68f
C335 w_611_305# p1g0 1.482f
C336 w_205_450# p2 1.014f
C337 w_569_n357# a_582_n389# 1.88f
C338 w_368_604# p3 1.014f
C339 w_678_68# a_691_36# 1.88f
C340 w_741_654# vdd 1.128f
C341 w_877_383# a_883_389# 2.444f
C342 b1 a_324_n46# 2.925f
C343 w_400_185# pocin 1.88f
C344 w_599_n75# a_579_n113# 1.014f
C345 w_258_17# vdd 1.128f
C346 w_642_625# p3p2p1g0 1.88f
C347 w_620_464# a_534_474# 3.59f
C348 w_877_383# a_825_350# 1.88f
C349 w_642_625# vdd 1.128f
C350 w_611_305# a_617_318# 1.41f
C351 w_400_185# a_380_153# 1.014f
C352 w_569_n357# a3 1.014f
C353 w_401_n240# vdd 1.128f
C354 w_400_323# p1g0 1.88f
C355 w_785_132# vdd 1.128f
C356 w_521_464# a_534_474# 2.45f
C357 w_879_518# a_884_498# 1.41f
C358 c2 s2 4.68f
C359 w_790_410# vdd 1.128f
C360 cin vdd 1.26f
C361 a1 b1 4.008f
C362 w_258_174# a_271_142# 1.88f
C363 g0 p1p0c0 0.18f
C364 w_329_n384# b3 1.17f
C365 w_538_625# vdd 1.128f
C366 p0 vdd 2.52f
C367 c2 a_815_n46# 1.845f
C368 a_612_n65# b1 2.674f
C369 w_400_28# a_324_88# 1.88f
C370 w_554_464# p1 1.014f
C371 w_329_n384# a3 1.128f
C372 w_367_n112# a_302_n114# 2.162f
C373 w_291_17# a_302_20# 1.014f
C374 w_439_167# vdd 1.41f
C375 w_400_28# b0 1.71f
C376 w_226_594# g2 2.268f
C377 g0 p1g0 1.01f
C378 w_238_456# g1 2.724f
C379 w_291_17# a_269_20# 1.88f
C380 w_506_301# a_453_311# 3.59f
C381 w_329_n250# p2 1.128f
C382 w_400_28# a0 1.014f
C383 w_434_604# vdd 1.128f
C384 w_417_462# a_397_472# 3.59f
C385 w_678_68# a_615_73# 1.014f
C386 a_206_556# g2 0.846f
C387 w_708_n70# vdd 1.128f
C388 w_599_n75# b1 1.128f
C389 a_304_190# vdd 1.89f
C390 w_258_174# p0 1.014f
C391 w_258_n117# a_269_n114# 1.014f
C392 w_726_513# vdd 1.88f
C393 w_797_280# cin 1.17f
C394 w_335_599# vdd 1.128f
C395 w_599_n75# a_612_n65# 2.82f
C396 w_566_n81# vdd 1.128f
C397 w_367_n112# b1 1.88f
C398 w_774_654# a_688_664# 3.59f
C399 a_239_604# g2 0.786f
C400 w_797_280# p0 1.128f
C401 w_401_n240# a_325_n180# 1.88f
C402 w_834_277# vdd 1.128f
C403 w_314_461# a_327_429# 1.88f
C404 a_600_239# gnd 1.616f
C405 w_367_n112# a1 1.17f
C406 w_587_464# vdd 1.128f
C407 w_401_n240# b2 1.71f
C408 w_193_588# vdd 1.128f
C409 w_711_68# g0 1.88f
C410 w_790_410# a_693_378# 1.014f
C411 w_258_312# a_271_280# 1.88f
C412 gnd 0 1.107555p **FLOATING
C413 g3 0 65.881004f **FLOATING
C414 vdd 0 0.797742p **FLOATING
C415 a_582_n389# 0 18.082f **FLOATING
C416 a_691_n378# 0 14.266f **FLOATING
C417 a_325_n314# 0 26.066f **FLOATING
C418 b3 0 90.43f **FLOATING
C419 a3 0 0.140213p **FLOATING
C420 a_615_n341# 0 44.863f **FLOATING
C421 a_582_n251# 0 18.082f **FLOATING
C422 a_325_n180# 0 26.066f **FLOATING
C423 b2 0 90.126f **FLOATING
C424 s3 0 21.761f **FLOATING
C425 a_831_n180# 0 26.066f **FLOATING
C426 a2 0 0.137957p **FLOATING
C427 c3 0 23.08f **FLOATING
C428 p3 0 0.410254p **FLOATING
C429 a_579_n113# 0 18.082f **FLOATING
C430 a_688_n102# 0 14.266f **FLOATING
C431 a_302_n114# 0 30.763f **FLOATING
C432 a_269_n114# 0 14.266f **FLOATING
C433 a_324_n46# 0 26.066f **FLOATING
C434 s2 0 20.539001f **FLOATING
C435 a_815_n46# 0 26.066f **FLOATING
C436 b1 0 93.114f **FLOATING
C437 a1 0 0.140495p **FLOATING
C438 a_612_n65# 0 44.863f **FLOATING
C439 c2 0 23.08f **FLOATING
C440 p2 0 0.53703p **FLOATING
C441 a_582_25# 0 18.082f **FLOATING
C442 a_691_36# 0 14.266f **FLOATING
C443 a_302_20# 0 30.763f **FLOATING
C444 a_269_20# 0 14.266f **FLOATING
C445 a_324_88# 0 26.066f **FLOATING
C446 b0 0 90.734f **FLOATING
C447 a0 0 0.144276p **FLOATING
C448 s1 0 20.539001f **FLOATING
C449 a_798_100# 0 26.066f **FLOATING
C450 a_615_73# 0 44.863f **FLOATING
C451 c1 0 23.08f **FLOATING
C452 a_445_140# 0 4.888f **FLOATING
C453 a_445_147# 0 20.28f **FLOATING
C454 p1 0 0.380473p **FLOATING
C455 pocin 0 28.03f **FLOATING
C456 a_271_142# 0 18.082f **FLOATING
C457 a_380_153# 0 14.266f **FLOATING
C458 a_496_232# 0 1.316f **FLOATING
C459 cin 0 85.827f **FLOATING
C460 p0 0 0.200305p **FLOATING
C461 s0 0 3.76f **FLOATING
C462 a_738_234# 0 26.066f **FLOATING
C463 a_304_190# 0 44.863f **FLOATING
C464 a_496_251# 0 1.316f **FLOATING
C465 p1p0c0 0 12.783999f **FLOATING
C466 a_617_278# 0 4.888f **FLOATING
C467 p1g0 0 18.06f **FLOATING
C468 a_600_239# 0 21.819f **FLOATING
C469 a_847_245# 0 14.266f **FLOATING
C470 a_771_282# 0 30.763f **FLOATING
C471 a_617_318# 0 2.585f **FLOATING
C472 g1 0 0.241318p **FLOATING
C473 a_453_311# 0 17.907999f **FLOATING
C474 a_271_280# 0 18.082f **FLOATING
C475 c4 0 4.324f **FLOATING
C476 p3p2p1p0c0 0 12.783999f **FLOATING
C477 a_380_291# 0 14.266f **FLOATING
C478 a_610_377# 0 1.128f **FLOATING
C479 g0 0 0.142494p **FLOATING
C480 a_304_328# 0 44.863f **FLOATING
C481 a_440_393# 0 1.316f **FLOATING
C482 a_610_395# 0 1.316f **FLOATING
C483 a_883_389# 0 4.888f **FLOATING
C484 p3p2p1g0 0 18.624f **FLOATING
C485 a_825_350# 0 23.605001f **FLOATING
C486 p2g1 0 12.22f **FLOATING
C487 a_610_414# 0 1.316f **FLOATING
C488 a_440_412# 0 1.316f **FLOATING
C489 a_731_417# 0 4.888f **FLOATING
C490 p2p1p0c0 0 18.624f **FLOATING
C491 a_883_429# 0 2.585f **FLOATING
C492 p3p2g1 0 30.286f **FLOATING
C493 a_693_378# 0 22.75f **FLOATING
C494 a_731_457# 0 2.585f **FLOATING
C495 p2p1g0 0 30.286f **FLOATING
C496 a_883_464# 0 2.35f **FLOATING
C497 p3g2 0 40.25f **FLOATING
C498 a_218_418# 0 18.082f **FLOATING
C499 a_534_474# 0 18.762999f **FLOATING
C500 a_397_472# 0 17.907999f **FLOATING
C501 a_327_429# 0 14.266f **FLOATING
C502 a_731_492# 0 2.35f **FLOATING
C503 g2 0 0.261375p **FLOATING
C504 a_884_498# 0 2.115f **FLOATING
C505 a_251_466# 0 44.863f **FLOATING
C506 a_424_535# 0 1.316f **FLOATING
C507 a_594_537# 0 1.316f **FLOATING
C508 a_797_547# 0 1.316f **FLOATING
C509 a_594_556# 0 1.316f **FLOATING
C510 a_424_554# 0 1.316f **FLOATING
C511 a_797_566# 0 1.316f **FLOATING
C512 a_594_575# 0 1.316f **FLOATING
C513 a_797_585# 0 1.316f **FLOATING
C514 a_797_604# 0 1.316f **FLOATING
C515 a_206_556# 0 18.082f **FLOATING
C516 a_315_567# 0 14.266f **FLOATING
C517 a_381_614# 0 17.907999f **FLOATING
C518 a_239_604# 0 44.863f **FLOATING
C519 a_518_635# 0 18.762999f **FLOATING
C520 a_688_664# 0 19.618f **FLOATING
