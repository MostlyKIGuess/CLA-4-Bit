* SPICE3 file created from cla.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Power Supply for the circuit
Vdd vdd gnd 'SUPPLY'


* Input Signals
* for testing
* Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
* Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 30n 60n)     
* Va1 a1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 10n 20n)    
* Vb1 b1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 30n 60n)    
* Va2 a2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 10n 20n)   
* Vb2 b2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 30n 60n)   
* Va3 a3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 10n 20n)   
* Vb3 b3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 30n 60n)   
* Vcin cin gnd DC 0         

* Input Signals for delay measurement

*  falling and rising
Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
Va1 a1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
Vb1 b1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
Va2 a2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Vb2 b2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Va3 a3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Vb3 b3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
Vcin cin gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)






* NGSPICE file created from testing.ext - technology: scmos

.option scale=90n

M1000 a_594_537# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1001 a_239_604# p3 g2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_329_n305# a_325_n314# p3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 a_218_418# p2 vdd w_205_450# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_825_350# g3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 a_600_239# p1p0c0 a_617_278# w_611_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 s1 p1 c1 w_818_n75# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 c1 a_445_147# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1008 p3p2p1g0 a_518_635# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1009 a_693_378# p2g1 a_731_417# w_725_411# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_564_n251# a2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1011 a_600_239# p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 a_594_n65# a1 b1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 gnd a_269_20# p0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 a_594_556# p2 a_594_537# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 a_445_147# g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1016 a_594_575# p1 a_594_556# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1017 p2g1 a_327_429# vdd w_347_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1018 a_440_412# p1 a_440_393# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_564_n389# a3 vdd w_551_n357# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1020 p1p0c0 a_453_311# vdd w_544_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1021 a3 b3 p3 w_329_n384# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 a_518_635# p3 vdd w_505_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a_731_457# p2p1p0c0 a_731_417# w_725_444# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1024 a_808_n381# p3 vdd w_795_n349# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1025 b2 a2 p2 w_368_n246# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1026 p3p2g1 a_381_614# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 p2p1p0c0 a_534_474# vdd w_658_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1028 a_610_395# p1 a_610_377# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1029 a_329_n171# a_325_n180# p2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 a_518_635# g0 a_594_575# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 s2 a_795_n247# a_873_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 vdd a0 a_324_88# w_400_28# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1033 a_594_n65# a_561_n113# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1034 vdd a_302_20# a_269_20# w_291_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 a_325_n180# b2 p2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 a_825_350# p3p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1037 a_304_190# a_271_142# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1038 a_847_245# a_771_282# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1039 a_884_498# p3g2 a_883_464# w_878_485# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 a_731_492# p2p1g0 a_731_457# w_725_479# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1041 a_673_n378# a_597_n341# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 a_597_n341# a_564_n389# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1043 a_315_567# a_239_604# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 g0 a_673_36# vdd w_693_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 p3g2 a_315_567# vdd w_335_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 vdd g3 a_884_498# w_879_518# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1047 a_825_350# p3p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 pocin a_380_153# vdd w_400_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 vdd a_269_20# p0 w_258_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 a_218_418# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1051 a_380_153# a_304_190# vdd w_367_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 b1 a1 a_302_n114# w_367_n112# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_825_350# p3p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1054 a_271_280# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1055 p3p2p1g0 a_518_635# vdd w_642_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_239_604# a_206_556# g2 w_226_594# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 a_304_190# a_271_142# cin w_291_180# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 c3 a_693_378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 g3 a_673_n378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 p2p1g0 a_397_472# vdd w_488_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_440_393# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_688_664# p0 vdd w_774_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 s2 p2 c2 w_815_n209# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1064 a_445_147# pocin gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 p2g1 a_327_429# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 a_600_239# p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1067 a_795_n247# p2 vdd w_782_n215# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_564_n251# a2 vdd w_551_n219# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_327_429# a_251_466# vdd w_314_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 a_688_664# cin vdd w_807_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1071 a_693_378# p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_251_466# p2 g1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 s1 c1 a_798_n113# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_798_n113# p1 vdd w_785_n81# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_325_n314# b3 p3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 a_738_234# p0 vdd w_725_266# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1077 a_673_36# a_597_73# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1078 a_564_25# a0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1079 p3p2g1 a_381_614# vdd w_472_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1080 a_597_n341# a_564_n389# b3 w_584_n351# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1081 a_206_556# p3 vdd w_193_588# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_424_535# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1083 g2 a_564_n251# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1084 g1 a_670_n102# vdd w_690_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1085 s3 p3 c3 w_828_n343# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_610_377# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1087 s0 a_847_245# vdd w_867_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1088 vdd a2 a_325_n180# w_401_n240# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_670_n102# a_594_n65# vdd w_657_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 c4 a_825_350# vdd w_942_382# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_670_n102# a_594_n65# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_424_554# p2 a_424_535# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 a_453_311# p0 vdd w_473_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1094 a_315_567# a_239_604# vdd w_302_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 p3p2p1p0c0 a_688_664# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_771_282# p0 cin w_758_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1097 s1 c1 p1 w_857_n67# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_271_142# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1099 a_534_474# cin vdd w_620_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_534_474# p0 vdd w_587_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_453_311# cin vdd w_506_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1102 a_271_280# p1 vdd w_258_312# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_561_n113# a1 vdd w_548_n81# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 a_381_614# g1 a_424_554# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_883_429# p3p2p1g0 a_883_389# w_877_416# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_693_378# p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 c1 a_445_147# vdd w_504_133# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_304_328# a_271_280# g0 w_291_318# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 a_825_350# p3g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1110 a_564_n389# a3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 s1 a_798_n113# a_876_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_688_664# p1 vdd w_741_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1113 a_797_604# p0 a_797_585# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 vdd a_269_n114# p1 w_258_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1115 p1g0 a_380_291# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_324_n46# b1 a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 a_327_429# a_251_466# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1118 a_693_378# p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 a_380_291# a_304_328# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1120 c2 a_600_239# vdd w_676_271# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 b3 a3 p3 w_368_n380# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1122 a1 b1 a_302_n114# w_328_n116# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 a_328_n37# a_324_n46# a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1124 a_328_97# a_324_88# a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 vdd a3 a_325_n314# w_401_n374# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1126 a_597_n341# a3 b3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 p1p0c0 a_453_311# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1128 a_324_88# b0 a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1129 a_688_664# cin a_797_604# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 vdd g2 a_731_492# w_726_513# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1131 a_883_464# p3p2g1 a_883_429# w_877_451# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_693_378# g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_304_328# p1 g0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1134 g2 a_564_n251# b2 w_584_n213# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1135 a_597_73# a_564_25# b0 w_584_63# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1136 a_597_73# a0 b0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1137 a_771_282# a_738_234# a_816_233# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1138 a_518_635# p1 vdd w_571_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_397_472# g0 vdd w_450_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_797_547# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_496_251# p0 a_496_232# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 a_847_245# a_771_282# vdd w_834_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_597_73# a_564_25# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1147 a_239_604# a_206_556# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1148 a_797_566# p2 a_797_547# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1149 a_453_311# cin a_496_251# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1150 a_453_311# p1 vdd w_440_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 gnd a3 a_325_n314# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1152 a_534_474# p1 vdd w_554_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_304_328# a_271_280# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1154 a_445_147# g0 a_445_140# w_439_134# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 a_797_585# p1 a_797_566# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 gnd a_302_n114# a_269_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_795_n247# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1158 gnd a_269_n114# p1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1159 g0 a_673_36# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1160 a_381_614# g1 vdd w_434_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 s2 c2 a_795_n247# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_561_n113# a1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1163 pocin a_380_153# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_380_153# a_304_190# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1165 a_688_664# p3 vdd w_675_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1166 s3 a_808_n381# a_886_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1167 a_673_n378# a_597_n341# vdd w_660_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 g2 a2 b2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 p1g0 a_380_291# vdd w_400_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1170 c2 a_600_239# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 g1 a_670_n102# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1172 a0 b0 a_302_20# w_328_18# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 a_380_291# a_304_328# vdd w_367_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_688_664# p2 vdd w_708_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1175 p2p1g0 a_397_472# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1176 gnd a2 a_325_n180# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 vdd pocin a_445_140# w_439_167# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1178 c3 a_693_378# vdd w_790_410# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_304_190# p0 cin Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1180 s3 c3 a_808_n381# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1181 a_251_466# a_218_418# g1 w_238_456# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1182 s3 c3 p3 w_867_n335# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 vdd a1 a_324_n46# w_400_n106# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1184 a_673_36# a_597_73# vdd w_660_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1185 a_397_472# g0 a_440_412# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 a_808_n381# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1187 a_798_n113# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_564_25# a0 vdd w_551_57# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 g3 a_673_n378# vdd w_693_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# p2 vdd w_384_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 vdd a_302_n114# a_269_n114# w_291_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1192 a_617_318# p1g0 a_617_278# w_611_305# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1193 a_771_282# cin p0 w_797_280# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 a_738_234# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1195 a_594_n65# a_561_n113# b1 w_581_n75# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_518_635# p2 vdd w_538_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 b0 a0 a_302_20# w_367_22# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_496_232# p1 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1199 a_397_472# p1 vdd w_417_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_206_556# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1201 p3p2p1p0c0 a_688_664# vdd w_845_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 a_610_414# p0 a_610_395# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_534_474# p2 vdd w_521_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_271_142# p0 vdd w_258_174# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1205 s0 a_847_245# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 vdd g1 a_617_318# w_611_340# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 c4 a_825_350# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1208 gnd a1 a_324_n46# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1209 gnd a0 a_324_88# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 gnd a_302_20# a_269_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1211 a_381_614# p2 vdd w_401_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1212 a2 b2 p2 w_329_n250# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 a_251_466# a_218_418# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 a_534_474# cin a_610_414# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1215 a_771_282# cin a_738_234# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 a_381_614# p3 vdd w_368_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1217 p3g2 a_315_567# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1218 a_600_239# g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1219 s2 c2 p2 w_854_n201# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 a_424_554# g1 0.013746f
C1 g3 p3p2g1 0.010274f
C2 a_594_537# gnd 0.412628f
C3 a_884_498# p3g2 3.63e-19
C4 g3 c2 0.005387f
C5 a_324_88# a0 0.060798f
C6 w_676_271# c2 0.016933f
C7 p1 vdd 0.796513f
C8 a_883_464# w_877_451# 0.01128f
C9 w_400_323# vdd 0.008451f
C10 a_795_n247# a_873_n248# 0.14502f
C11 w_367_22# a_302_20# 0.015055f
C12 w_367_n112# a1 0.028748f
C13 w_328_n116# b1 0.027716f
C14 vdd w_521_464# 0.008451f
C15 p2p1g0 gnd 0.210726f
C16 a_883_464# p3p2p1g0 0.016011f
C17 p0 w_584_63# 0.00465f
C18 a_218_418# gnd 0.208267f
C19 w_367_185# vdd 0.008465f
C20 a_884_498# vdd 0.41238f
C21 a_304_328# vdd 0.017291f
C22 w_725_266# vdd 0.008698f
C23 a_600_239# p1p0c0 0.211061f
C24 p3g2 p3p2p1g0 0.001431f
C25 p2p1g0 a_397_472# 0.060798f
C26 p1 a_798_n113# 0.060798f
C27 a_847_245# gnd 0.248155f
C28 w_818_n75# c1 0.015306f
C29 w_587_464# g2 0.00583f
C30 a_327_429# p2g1 0.060798f
C31 a_564_n389# vdd 0.439906f
C32 a_693_378# vdd 0.001532f
C33 vdd w_877_451# 0.010901f
C34 g2 g1 1.67738f
C35 a_688_664# a_797_604# 0.41238f
C36 w_238_456# g1 0.021496f
C37 vdd a_453_311# 1.32165f
C38 w_314_461# g2 0.005799f
C39 p1 a_797_566# 0.013746f
C40 cin a_797_585# 2.05e-21
C41 a_886_n382# s3 0.20619f
C42 p0 a_738_234# 0.060798f
C43 vdd p3p2p1g0 0.4601f
C44 a2 a_564_n251# 0.060825f
C45 b2 a_329_n171# 0.001802f
C46 a_884_498# w_878_485# 0.01128f
C47 g0 w_658_464# 0.002547f
C48 p3 a_315_567# 0.001362f
C49 p2 a_381_614# 0.005763f
C50 w_807_654# vdd 0.008451f
C51 w_551_n219# a_564_n251# 0.013216f
C52 a_731_492# vdd 0.41238f
C53 a_731_457# w_725_444# 0.009864f
C54 gnd a_670_n102# 0.248155f
C55 c2 s1 0.002762f
C56 p3p2p1g0 w_878_485# 0.011197f
C57 vdd b0 0.019072f
C58 w_258_n117# vdd 0.008451f
C59 cin w_400_185# 0.00869f
C60 w_828_n343# c3 0.016729f
C61 w_401_n240# vdd 0.026104f
C62 w_329_n250# a2 0.007896f
C63 cin c3 5.08e-19
C64 g0 a_440_412# 0.014522f
C65 w_795_n349# p3 0.028034f
C66 a_876_n114# a_798_n113# 0.14502f
C67 g2 w_488_462# 0.005809f
C68 p1 p2 2.60374f
C69 p0 p3 0.002227f
C70 p3p2p1p0c0 w_879_518# 0.015324f
C71 w_434_604# vdd 0.008451f
C72 g3 g2 0.005441f
C73 a_251_466# g1 0.770057f
C74 a_251_466# w_314_461# 0.026907f
C75 p2 w_521_464# 0.026794f
C76 p0 g0 0.074894f
C77 p1 a_518_635# 0.005763f
C78 w_611_340# a_617_318# 0.009864f
C79 cin a_688_664# 0.059029f
C80 w_329_n384# a3 0.007896f
C81 w_611_305# p1p0c0 1.04e-20
C82 a1 vdd 0.230834f
C83 w_797_280# c3 0.012687f
C84 g2 b3 3.99e-19
C85 vdd a_380_153# 0.443425f
C86 a_564_25# b0 0.00288f
C87 p0 a_597_73# 0.007562f
C88 g0 a_445_147# 0.216537f
C89 s3 c3 0.692464f
C90 p2g1 w_347_461# 0.013223f
C91 g0 a_610_377# 0.002334f
C92 w_867_n335# s3 0.007992f
C93 p3 a_808_n381# 0.060798f
C94 p3g2 g1 0.023512f
C95 g2 w_193_588# 0.009535f
C96 a_825_350# p3p2p1p0c0 0.217915f
C97 p1 w_258_312# 0.028034f
C98 a_883_389# p3p2p1g0 0.004158f
C99 c3 gnd 0.42764f
C100 c3 a_795_n247# 4.01e-19
C101 b1 a_561_n113# 0.00343f
C102 p1 w_417_462# 0.026996f
C103 w_587_464# vdd 0.008451f
C104 p2 p3p2p1g0 0.010267f
C105 w_258_17# vdd 0.008451f
C106 p2p1p0c0 a_731_417# 0.004158f
C107 g0 p1p0c0 0.010775f
C108 cin a_771_282# 0.68509f
C109 a_534_474# a_610_414# 0.41238f
C110 cin a_797_547# 2.48e-20
C111 p2g1 a_731_417# 0.019622f
C112 w_314_461# vdd 0.012946f
C113 w_690_n70# a_670_n102# 0.026907f
C114 a_518_635# p3p2p1g0 0.060798f
C115 vdd g1 0.886292f
C116 a_688_664# gnd 0.042086f
C117 p3 w_505_625# 0.026794f
C118 w_400_n106# vdd 0.026082f
C119 p0 p2p1g0 0.009782f
C120 gnd c1 0.261394f
C121 cin a_534_474# 0.060518f
C122 p1 p2g1 0.03968f
C123 w_797_280# a_771_282# 0.007992f
C124 c4 gnd 0.302435f
C125 w_401_n240# p2 0.003504f
C126 a3 b3 0.535308f
C127 p0 a_328_97# 3.98e-19
C128 a_315_567# w_302_599# 0.013216f
C129 a_206_556# w_226_594# 0.026794f
C130 a_564_n389# a_597_n341# 0.003752f
C131 w_548_n81# a_561_n113# 0.013216f
C132 a_329_n305# b3 0.001802f
C133 w_400_185# pocin 0.013216f
C134 w_611_272# p1g0 0.001158f
C135 a_797_547# gnd 0.41238f
C136 g3 p3g2 0.013767f
C137 gnd a_771_282# 0.190422f
C138 p2p1p0c0 a_693_378# 0.040556f
C139 b0 a0 0.539271f
C140 a_693_378# p2g1 0.244568f
C141 w_367_323# vdd 0.008493f
C142 w_400_28# a_324_88# 0.013216f
C143 a_795_n247# s2 0.286223f
C144 w_328_18# a_302_20# 0.007992f
C145 w_328_n116# a1 0.007896f
C146 p2 a_594_556# 0.023173f
C147 vdd w_488_462# 0.008451f
C148 a_883_464# p3p2g1 3.63e-19
C149 a_534_474# gnd 0.042086f
C150 w_291_180# vdd 6.13e-19
C151 g3 vdd 0.487338f
C152 a_617_278# p1g0 0.004158f
C153 w_676_271# vdd 0.008511f
C154 gnd a_325_n180# 0.206673f
C155 p3g2 p3p2g1 0.633236f
C156 vdd b3 0.016782f
C157 p1 a_561_n113# 0.002494f
C158 w_554_464# g2 0.0039f
C159 gnd a_302_20# 0.190422f
C160 a_673_n378# vdd 0.441438f
C161 vdd w_790_410# 0.008495f
C162 w_782_n215# a_795_n247# 0.013216f
C163 w_205_450# g1 0.013044f
C164 w_238_456# g2 0.001868f
C165 p0 a_797_585# 0.013746f
C166 vdd p1g0 0.451968f
C167 p1 a_594_575# 0.031835f
C168 cin a_797_604# 0.013759f
C169 a_886_n382# a_808_n381# 0.14502f
C170 vdd p3p2g1 0.454731f
C171 vdd w_193_588# 0.0086f
C172 c2 vdd 0.442422f
C173 b2 a_325_n180# 0.02927f
C174 p3 w_368_n380# 0.015055f
C175 cin w_726_513# 0.002754f
C176 w_774_654# vdd 0.008451f
C177 p2 g1 0.146262f
C178 p3 a_381_614# 0.003255f
C179 a_816_233# a_738_234# 0.14502f
C180 a_269_20# a_302_20# 0.060798f
C181 a_324_88# a_328_97# 0.14502f
C182 p2p1p0c0 w_725_411# 0.001174f
C183 a_269_n114# gnd 0.248155f
C184 w_725_266# a_738_234# 0.013216f
C185 p0 w_611_340# 1.24e-20
C186 p2g1 w_725_411# 0.049155f
C187 a_884_498# w_879_518# 0.009864f
C188 c2 a_798_n113# 0.003242f
C189 p3p2g1 w_878_485# 6.13e-19
C190 w_693_68# vdd 0.008451f
C191 w_584_63# b0 0.008938f
C192 cin a_610_414# 0.013746f
C193 p0 c3 1.47e-20
C194 a_731_492# w_725_479# 0.01128f
C195 g1 w_417_462# 2.78e-19
C196 g2 w_450_462# 0.005809f
C197 p1 p3 0.040972f
C198 p3p2p1g0 w_879_518# 0.011197f
C199 a_251_466# w_238_456# 0.019526f
C200 w_401_604# vdd 0.008451f
C201 a_251_466# g2 0.005106f
C202 p2p1g0 w_620_464# 9.19e-21
C203 gnd a_206_556# 0.20619f
C204 p1 g0 0.060865f
C205 p0 a_688_664# 0.005763f
C206 a_594_n65# vdd 0.013824f
C207 g2 a3 0.009821f
C208 a_534_474# w_658_464# 0.027163f
C209 g0 w_400_323# 0.011443f
C210 g3 p2 0.022389f
C211 g1 w_384_462# 0.011399f
C212 p2 a_440_393# 0.013746f
C213 a_798_n113# s1 0.286223f
C214 a_808_n381# c3 0.017003f
C215 p0 c1 0.015446f
C216 p2g1 g1 0.007851f
C217 g0 a_304_328# 0.753587f
C218 cin w_797_280# 0.027729f
C219 w_828_n343# s3 0.015055f
C220 a_600_239# g1 1.39e-20
C221 a_445_147# c1 0.060798f
C222 a_825_350# p3p2p1g0 0.040556f
C223 a_324_n46# a_328_n37# 0.14502f
C224 a_269_n114# a_302_n114# 0.060798f
C225 a1 a_561_n113# 0.060856f
C226 w_554_464# vdd 0.008451f
C227 a_302_n114# a_328_n37# 0.20619f
C228 p2 p3p2g1 0.017215f
C229 p3 p3p2p1g0 0.010267f
C230 p2 c2 0.026943f
C231 w_504_133# vdd 0.008451f
C232 p0 a_771_282# 0.413834f
C233 a_594_575# a_594_556# 0.41238f
C234 w_238_456# vdd 6.13e-19
C235 vdd g2 0.07536f
C236 cin gnd 0.067929f
C237 g0 p3p2p1g0 0.001581f
C238 a_518_635# p3p2g1 0.041586f
C239 a_688_664# p3p2p1p0c0 0.060798f
C240 w_367_n112# vdd 6.13e-19
C241 p1 p2p1g0 0.016236f
C242 p0 a_534_474# 0.005763f
C243 w_758_272# a_771_282# 0.015055f
C244 a_380_291# gnd 0.248155f
C245 p2p1g0 w_521_464# 1.11e-19
C246 w_291_318# a_271_280# 0.026794f
C247 a_597_n341# b3 0.756931f
C248 p0 a_302_20# 0.003749f
C249 a_673_n378# a_597_n341# 0.060798f
C250 a_325_n314# b3 0.02927f
C251 p3p2p1g0 w_642_625# 0.013284f
C252 p2p1p0c0 a_731_457# 4.37e-21
C253 p2p1g0 a_693_378# 0.001345f
C254 b0 a_597_73# 0.756776f
C255 w_676_271# a_600_239# 0.027289f
C256 w_611_272# a_617_278# 0.017071f
C257 p2 w_401_604# 0.026996f
C258 gnd a_795_n247# 0.206673f
C259 w_291_318# vdd 6.13e-19
C260 w_291_17# a_302_20# 0.027261f
C261 w_400_28# b0 0.015139f
C262 p2 a_424_554# 0.023081f
C263 p3 a_594_556# 0.016756f
C264 vdd w_450_462# 0.008451f
C265 p1 w_857_n67# 0.007896f
C266 a_397_472# gnd 0.042086f
C267 a_251_466# vdd 0.019451f
C268 w_258_174# vdd 0.009216f
C269 w_611_305# g1 0.002086f
C270 a_600_239# p1g0 0.040556f
C271 cin pocin 0.002387f
C272 gnd b2 0.039557f
C273 vdd a3 0.209306f
C274 p2p1g0 a_731_492# 3.63e-19
C275 p1 a_670_n102# 0.002494f
C276 a_600_239# c2 0.060798f
C277 gnd a_269_20# 0.248155f
C278 a_883_464# vdd 0.014511f
C279 a_445_140# pocin 0.185571f
C280 w_854_n201# c2 0.027735f
C281 w_205_450# g2 0.001868f
C282 vdd a_271_280# 0.455487f
C283 a_239_604# g2 0.75303f
C284 p1 a_797_585# 0.013746f
C285 p0 a_797_604# 0.013746f
C286 vdd p3g2 0.447846f
C287 a2 a_325_n180# 0.060798f
C288 p3 w_329_n384# 0.007992f
C289 p2 g2 0.077377f
C290 p3 g1 0.658617f
C291 w_741_654# vdd 0.008451f
C292 a_424_535# a_424_554# 0.41238f
C293 a_594_537# a_594_556# 0.41238f
C294 w_584_n213# b2 0.008451f
C295 a_324_88# a_302_20# 0.286223f
C296 a_731_457# w_725_479# 0.009864f
C297 p2p1p0c0 w_725_444# 0.036782f
C298 g0 g1 6.14e-19
C299 b0 a_328_97# 0.001802f
C300 w_693_68# a_673_36# 0.026907f
C301 a_883_464# w_878_485# 0.009864f
C302 a_324_n46# gnd 0.206673f
C303 cin w_506_301# 0.026794f
C304 gnd pocin 0.386422f
C305 g3 w_879_518# 0.036563f
C306 gnd a_302_n114# 0.190422f
C307 p3g2 w_878_485# 0.036563f
C308 w_660_68# vdd 0.02492f
C309 p3p2g1 a_594_575# 7.98e-19
C310 p3g2 a_797_566# 0.004452f
C311 p0 a_610_414# 0.019134f
C312 a_564_n389# w_584_n351# 0.026794f
C313 a_673_n378# w_660_n346# 0.013216f
C314 vdd a_798_n113# 0.442386f
C315 c2 a_738_234# 0.003282f
C316 g2 w_417_462# 0.005809f
C317 a_269_n114# w_291_n117# 0.013216f
C318 p3p2g1 w_879_518# 4.09e-19
C319 w_368_604# vdd 0.008451f
C320 p2p1g0 w_587_464# 8.56e-21
C321 w_611_305# p1g0 0.036784f
C322 g3 a_825_350# 0.001813f
C323 w_544_301# p1p0c0 0.013229f
C324 gnd a_315_567# 0.248155f
C325 p1 a_688_664# 0.004034f
C326 p0 cin 0.257529f
C327 g2 a_597_n341# 0.013288f
C328 a_564_25# vdd 0.439891f
C329 a_534_474# w_620_464# 0.027639f
C330 g0 w_367_323# 0.011382f
C331 vdd s0 0.439883f
C332 a_251_466# p2 0.001371f
C333 g2 w_384_462# 0.005809f
C334 p2p1p0c0 g2 0.065766f
C335 p1 c1 0.024407f
C336 p3 b3 0.685112f
C337 a_693_378# c3 0.060798f
C338 p2g1 g2 0.00516f
C339 a_218_418# g1 0.012164f
C340 g0 g3 0.00202f
C341 p0 w_797_280# 0.007968f
C342 cin w_758_272# 0.013523f
C343 g0 a_440_393# 7.76e-19
C344 g2 a_564_n251# 0.003752f
C345 a_445_147# a_445_140# 0.453641f
C346 a_825_350# p3p2g1 0.001345f
C347 a_440_412# gnd 1.91e-19
C348 a_594_n65# a_561_n113# 0.003752f
C349 b1 a_328_n37# 0.001802f
C350 a_324_n46# a_302_n114# 0.286223f
C351 p3 w_193_588# 0.028034f
C352 p3 p3p2g1 0.017448f
C353 p2 p3g2 0.026294f
C354 a_397_472# a_440_412# 0.41238f
C355 cin p1p0c0 0.013387f
C356 g0 p1g0 0.015977f
C357 w_205_450# vdd 0.0086f
C358 a_688_664# p3p2p1g0 0.00431f
C359 g0 p3p2g1 0.015172f
C360 vdd a_239_604# 0.024911f
C361 a_518_635# p3g2 8.1e-19
C362 p0 gnd 0.898603f
C363 cin a_304_190# 0.747651f
C364 c3 a_876_n114# 6.44e-19
C365 w_328_n116# vdd 0.001288f
C366 a_688_664# w_807_654# 0.027639f
C367 a_816_233# a_771_282# 0.20619f
C368 p2 vdd 0.774066f
C369 gnd a_445_147# 0.576829f
C370 g3 w_834_277# 0.016049f
C371 p1 a_534_474# 0.015195f
C372 a_808_n381# s3 0.286223f
C373 a_610_377# gnd 0.41238f
C374 p2p1g0 w_488_462# 0.013216f
C375 a_518_635# vdd 1.76176f
C376 w_845_654# vdd 0.008451f
C377 w_258_312# a_271_280# 0.013216f
C378 a_534_474# w_521_464# 0.017642f
C379 g1 a_670_n102# 0.060798f
C380 p2 w_368_n246# 0.018553f
C381 a_597_n341# a3 0.001371f
C382 a_808_n381# gnd 0.206673f
C383 p0 a_269_20# 0.06476f
C384 a_325_n314# a3 0.060798f
C385 g0 w_693_68# 0.01325f
C386 vdd a0 0.236105f
C387 w_400_185# a_380_153# 0.026907f
C388 a_876_n114# c1 0.001856f
C389 p3p2p1p0c0 w_877_383# 0.053825f
C390 a_325_n314# a_329_n305# 0.14502f
C391 w_551_57# vdd 0.0086f
C392 g3 a_847_245# 0.015251f
C393 gnd p1p0c0 0.207724f
C394 w_834_277# c2 8.35e-21
C395 w_611_272# a_600_239# 0.013329f
C396 p3p2p1p0c0 gnd 0.216485f
C397 w_258_312# vdd 0.028134f
C398 a_304_190# gnd 0.701773f
C399 w_291_17# a_269_20# 0.013216f
C400 w_367_22# b0 0.01395f
C401 c2 a_873_n248# 0.001866f
C402 p2 a_797_566# 0.013746f
C403 p3 a_424_554# 0.025115f
C404 vdd w_417_462# 0.008451f
C405 p1 w_818_n75# 0.028748f
C406 a_327_429# gnd 0.248155f
C407 w_867_277# vdd 0.008451f
C408 p1 a_269_n114# 0.06333f
C409 w_611_340# g1 0.039692f
C410 cin a_271_142# 0.001372f
C411 gnd a2 1.55938f
C412 p0 pocin 5.46e-21
C413 vdd a_597_n341# 0.011744f
C414 p1 a_328_n37# 6.43e-21
C415 a_600_239# a_617_278# 0.453641f
C416 a_564_25# a0 0.060867f
C417 a_325_n314# vdd 0.442574f
C418 vdd w_384_462# 0.008451f
C419 gnd a_324_88# 0.206673f
C420 p2p1p0c0 vdd 0.439883f
C421 a_445_147# pocin 1.39e-20
C422 p2g1 vdd 0.439883f
C423 w_815_n209# c2 0.01623f
C424 w_551_57# a_564_25# 0.013216f
C425 vdd a_564_n251# 0.455188f
C426 a2 b2 0.531092f
C427 a_600_239# vdd 0.001532f
C428 cin w_620_464# 0.026794f
C429 p2 w_205_450# 0.028034f
C430 p3 g2 0.017978f
C431 w_708_654# vdd 0.008451f
C432 g0 w_504_133# 0.011197f
C433 vdd a_673_36# 0.441647f
C434 w_401_n240# a_325_n180# 0.013216f
C435 b0 a_302_20# 0.685117f
C436 g0 g2 0.017633f
C437 w_660_68# a_673_36# 0.013216f
C438 w_867_277# s0 0.013216f
C439 b1 gnd 0.03874f
C440 gnd a_271_142# 0.20619f
C441 p1 w_657_n70# 0.002922f
C442 g1 c1 0.008592f
C443 a_518_635# p2 0.004034f
C444 w_584_63# vdd 2.04e-19
C445 w_335_599# p3g2 0.013277f
C446 w_584_n351# b3 0.008451f
C447 p3p2g1 a_797_585# 0.049949f
C448 p3p2p1g0 a_797_604# 0.043431f
C449 p3g2 a_594_575# 0.042464f
C450 a_564_n389# w_551_n357# 0.013216f
C451 vdd a_561_n113# 0.439891f
C452 a_269_n114# w_258_n117# 0.026907f
C453 w_335_599# vdd 0.008451f
C454 w_291_n117# a_302_n114# 0.027261f
C455 g3 c3 0.073145f
C456 p2p1g0 w_554_464# 8.56e-21
C457 w_544_301# a_453_311# 0.027163f
C458 w_857_n67# s1 0.007992f
C459 gnd a_381_614# 0.042086f
C460 p1 cin 0.034484f
C461 a_534_474# w_587_464# 0.027639f
C462 g0 w_291_318# 0.008451f
C463 a_731_492# w_726_513# 0.009864f
C464 vdd a_738_234# 0.439891f
C465 w_611_305# a_617_278# 0.008113f
C466 w_551_57# a0 0.028093f
C467 a_424_535# p2 0.023137f
C468 g0 w_450_462# 0.026794f
C469 a_564_25# w_584_63# 0.026794f
C470 p2p1g0 g2 0.005084f
C471 cin a_816_233# 0.002154f
C472 vdd w_879_518# 0.013167f
C473 p0 a_445_147# 2.69e-20
C474 a_218_418# g2 0.002036f
C475 p3 a3 0.413834f
C476 a_218_418# w_238_456# 0.026794f
C477 c3 w_790_410# 0.013216f
C478 p0 a_610_377# 6.84e-20
C479 cin w_367_185# 0.00869f
C480 p2 w_384_462# 0.026794f
C481 w_660_n346# vdd 0.008611f
C482 p0 w_758_272# 0.028748f
C483 b1 a_324_n46# 0.02927f
C484 p3 a_329_n305# 0.20619f
C485 w_400_323# a_380_291# 0.026907f
C486 w_795_n349# a_808_n381# 0.013216f
C487 p2 p2g1 0.004909f
C488 a_825_350# p3g2 0.001345f
C489 a_594_n65# a_670_n102# 0.060798f
C490 b1 a_302_n114# 0.685112f
C491 c2 c3 0.026004f
C492 g3 c1 0.003696f
C493 w_439_167# vdd 0.0112f
C494 p2 a_564_n251# 0.002692f
C495 p3 p3g2 0.026608f
C496 a_304_328# a_380_291# 0.060798f
C497 p1 w_571_625# 0.026996f
C498 g0 a_271_280# 0.001372f
C499 cin a_453_311# 0.069062f
C500 w_708_654# p2 0.026794f
C501 p1 gnd 0.59676f
C502 cin p3p2p1g0 0.02473f
C503 g0 p3g2 0.0027f
C504 cin a_496_251# 0.014005f
C505 p0 a_304_190# 0.001371f
C506 a_825_350# vdd 0.011869f
C507 w_854_n201# p2 0.007896f
C508 cin w_807_654# 0.026794f
C509 a_688_664# w_774_654# 0.027639f
C510 p3 vdd 0.984731f
C511 g3 a_771_282# 2.33e-19
C512 p1 a_397_472# 0.017711f
C513 c2 c1 0.013027f
C514 a_304_328# gnd 0.588368f
C515 g0 vdd 0.632781f
C516 p2g1 w_417_462# 8.35e-22
C517 a_883_429# w_877_416# 0.009864f
C518 p2 w_329_n250# 0.011491f
C519 w_581_n75# b1 0.009938f
C520 c3 s1 0.003481f
C521 a_251_466# a_218_418# 0.003752f
C522 p0 a_324_88# 0.0179f
C523 a_564_n389# gnd 0.20619f
C524 a_693_378# gnd 1.08291f
C525 a_883_429# p3p2p1p0c0 0.005194f
C526 vdd a_597_73# 0.015633f
C527 p3p2p1p0c0 w_877_416# 0.018361f
C528 p3p2p1g0 w_877_383# 0.001142f
C529 gnd a_453_311# 0.042086f
C530 w_400_28# vdd 0.023245f
C531 w_660_68# a_597_73# 0.026907f
C532 c2 a_771_282# 0.020436f
C533 p2g1 w_384_462# 1.09e-20
C534 p3p2p1g0 gnd 0.232346f
C535 p2p1p0c0 p2g1 0.008706f
C536 p3 w_368_604# 0.026794f
C537 c2 s2 0.686118f
C538 w_328_18# b0 0.027757f
C539 c1 s1 0.686034f
C540 p1 w_785_n81# 0.028309f
C541 vdd w_642_625# 0.008451f
C542 a_518_635# a_594_575# 0.41238f
C543 p1 a_324_n46# 0.008083f
C544 w_834_277# vdd 0.008512f
C545 p0 a_271_142# 0.060798f
C546 cin a_380_153# 0.003392f
C547 p1 a_302_n114# 0.007287f
C548 gnd b0 0.045026f
C549 a_564_25# a_597_73# 0.003752f
C550 p2p1g0 vdd 0.439883f
C551 p1 w_690_n70# 0.002922f
C552 a_218_418# vdd 0.439891f
C553 a_825_350# a_883_389# 0.453641f
C554 a_847_245# vdd 0.441416f
C555 p3 a_239_604# 0.002112f
C556 w_675_654# vdd 0.008451f
C557 g0 w_439_134# 0.051057f
C558 w_551_n219# a2 0.028079f
C559 w_401_n240# b2 0.015139f
C560 w_815_n209# vdd 4.8e-19
C561 c2 w_818_n75# 0.019549f
C562 cin g1 0.016729f
C563 p3 p2 0.395341f
C564 a1 gnd 1.83674f
C565 p0 w_473_301# 0.026996f
C566 w_504_133# c1 0.013242f
C567 gnd a_380_153# 0.248155f
C568 a_304_190# a_271_142# 0.003752f
C569 p1 w_581_n75# 0.002922f
C570 g0 p2 0.045639f
C571 a_518_635# p3 0.002444f
C572 w_660_n346# a_597_n341# 0.026907f
C573 g0 a_518_635# 0.06069f
C574 p3p2g1 a_797_604# 0.003102f
C575 p3g2 a_797_585# 0.054573f
C576 p1 a_440_412# 0.013746f
C577 a_847_245# s0 0.060798f
C578 vdd a_670_n102# 0.441416f
C579 vdd w_302_599# 0.016007f
C580 g1 a_617_318# 0.010567f
C581 w_506_301# a_453_311# 0.027639f
C582 w_544_301# p1g0 0.004305f
C583 gnd g1 0.512437f
C584 p1 p0 0.069366f
C585 w_818_n75# s1 0.015055f
C586 a_206_556# w_193_588# 0.013216f
C587 a_597_73# a0 0.001371f
C588 a_534_474# w_554_464# 0.027639f
C589 p1 w_440_301# 0.026794f
C590 a_424_535# p3 0.013746f
C591 a_594_537# p2 0.020283f
C592 w_400_28# a0 0.028034f
C593 a_397_472# g1 0.007928f
C594 a_534_474# g2 0.009442f
C595 a_327_429# w_347_461# 0.026907f
C596 a_218_418# w_205_450# 0.013216f
C597 a_518_635# w_642_625# 0.027163f
C598 p1 a_610_377# 0.013746f
C599 cin w_291_180# 0.008451f
C600 p0 w_725_266# 0.028034f
C601 a1 a_324_n46# 0.060798f
C602 p3 a_325_n314# 0.286223f
C603 p2 p2p1g0 0.001781f
C604 w_258_17# a_269_20# 0.026907f
C605 w_367_323# a_380_291# 0.013216f
C606 g1 b2 7.83e-19
C607 w_611_340# vdd 0.066855f
C608 a1 a_302_n114# 0.413834f
C609 p2 a_218_418# 0.061185f
C610 a_380_153# pocin 0.060798f
C611 g0 p2p1p0c0 0.073898f
C612 p0 a_693_378# 6.43e-21
C613 p2 a_329_n171# 0.20619f
C614 w_400_185# vdd 0.02411f
C615 g0 p2g1 0.004954f
C616 a_797_585# a_797_566# 0.41238f
C617 p0 a_453_311# 0.005763f
C618 cin p1g0 0.012177f
C619 w_440_301# a_453_311# 0.017642f
C620 cin p3p2g1 0.004802f
C621 p0 p3p2p1g0 0.013325f
C622 p0 a_496_251# 0.013746f
C623 cin c2 0.003312f
C624 w_815_n209# p2 0.028748f
C625 c3 vdd 0.446488f
C626 g0 a_673_36# 0.060812f
C627 a_688_664# w_741_654# 0.027639f
C628 w_472_604# a_381_614# 0.027163f
C629 a_380_291# p1g0 0.060798f
C630 a_884_498# p3p2p1p0c0 0.005507f
C631 g3 gnd 0.253819f
C632 a_440_393# gnd 0.41811f
C633 w_367_185# a_304_190# 0.026907f
C634 a_673_36# a_597_73# 0.060798f
C635 w_797_280# c2 0.003455f
C636 a_688_664# vdd 2.20188f
C637 a_397_472# w_488_462# 0.027163f
C638 a_883_429# w_877_451# 0.009864f
C639 gnd b3 0.035921f
C640 w_400_n106# a_324_n46# 0.013216f
C641 w_657_n70# a_594_n65# 0.026907f
C642 c3 a_798_n113# 0.001329f
C643 p0 b0 0.023585f
C644 a_673_n378# gnd 0.248155f
C645 a_883_429# p3p2p1g0 0.00801f
C646 a_239_604# w_302_599# 0.026907f
C647 g2 w_226_594# 0.018971f
C648 vdd c1 0.444335f
C649 a_453_311# p1p0c0 0.060798f
C650 p3p2p1g0 w_877_416# 0.03763f
C651 p3p2p1p0c0 w_877_451# 0.018013f
C652 p1g0 a_617_318# 4.37e-21
C653 w_690_n70# g1 0.01323f
C654 gnd p1g0 0.207724f
C655 w_367_22# vdd 6.13e-19
C656 c4 vdd 0.439883f
C657 a_797_547# p3g2 0.001272f
C658 w_867_277# a_847_245# 0.026907f
C659 p2p1g0 p2p1p0c0 0.057637f
C660 w_584_63# a_597_73# 0.019526f
C661 p3p2p1g0 p3p2p1p0c0 0.003212f
C662 p3p2g1 gnd 0.234908f
C663 p2p1g0 p2g1 0.005273f
C664 c2 gnd 0.219293f
C665 c3 s0 0.003003f
C666 c2 a_795_n247# 0.017003f
C667 w_726_513# g2 0.036563f
C668 p3 a_594_575# 2.95e-20
C669 vdd w_942_382# 0.00851f
C670 vdd w_604_625# 0.008451f
C671 c1 a_798_n113# 0.016996f
C672 g2 a_206_556# 0.008991f
C673 g0 a_594_575# 0.013746f
C674 vdd a_771_282# 0.019283f
C675 p1 b1 0.022716f
C676 cin a_496_232# 0.024151f
C677 a_534_474# vdd 1.76176f
C678 vdd a_325_n180# 0.443244f
C679 p0 w_587_464# 0.026996f
C680 g0 w_439_167# 4.29e-19
C681 vdd a_302_20# 0.019283f
C682 p0 w_258_17# 0.013216f
C683 w_401_n240# a2 0.028034f
C684 a_797_547# a_797_566# 0.41238f
C685 w_782_n215# vdd 0.019776f
C686 b0 a_324_88# 0.02927f
C687 p0 g1 0.031532f
C688 cin g2 0.005207f
C689 p2p1g0 w_725_479# 0.036563f
C690 a_594_n65# gnd 0.701773f
C691 gnd a_496_232# 0.41238f
C692 a_304_190# a_380_153# 0.060798f
C693 p1 w_548_n81# 0.002922f
C694 a_688_664# p2 0.004034f
C695 g0 p3 0.057959f
C696 w_818_n75# vdd 8.63e-20
C697 a_688_664# w_845_654# 0.027163f
C698 w_401_n374# b3 0.015139f
C699 w_551_n357# a3 0.02808f
C700 w_584_n351# a_597_n341# 0.019526f
C701 a_269_n114# vdd 0.441416f
C702 vdd w_226_594# 6.13e-19
C703 g1 p1p0c0 0.002848f
C704 w_238_456# gnd 0.003687f
C705 w_473_301# a_453_311# 0.027639f
C706 a_440_393# a_440_412# 0.41238f
C707 w_867_277# c3 3.18e-20
C708 a_610_395# a_610_414# 0.41238f
C709 w_506_301# p1g0 0.004305f
C710 gnd g2 0.865158f
C711 a_797_547# p2 0.013746f
C712 a_594_537# p3 0.013776f
C713 w_367_22# a0 0.028748f
C714 w_726_513# vdd 0.013119f
C715 a_693_378# a_731_417# 0.453641f
C716 a_327_429# g1 0.009049f
C717 p2 s2 0.413834f
C718 a_327_429# w_314_461# 0.013216f
C719 a_397_472# g2 0.00724f
C720 a_518_635# w_604_625# 0.027639f
C721 p1 a_304_328# 0.04464f
C722 a1 b1 0.614689f
C723 w_551_n357# vdd 0.008823f
C724 vdd a_206_556# 0.439891f
C725 g2 b2 0.764942f
C726 g1 a2 0.011016f
C727 w_544_301# vdd 0.008451f
C728 p2 a_534_474# 0.002444f
C729 w_657_n70# vdd 0.008534f
C730 g0 p2p1g0 0.001609f
C731 p2 a_325_n180# 0.288532f
C732 w_584_n213# g2 0.019526f
C733 w_854_n201# c3 5.29e-20
C734 p0 p1g0 7.17e-19
C735 p1 a_453_311# 0.002444f
C736 w_675_654# p3 0.026794f
C737 w_440_301# p1g0 0.004305f
C738 cin p3g2 0.004802f
C739 p1 p3p2p1g0 0.010267f
C740 p0 p3p2g1 0.012004f
C741 p0 c2 0.020959f
C742 w_782_n215# p2 0.028034f
C743 a_688_664# w_708_654# 0.027639f
C744 p0 w_774_654# 0.026996f
C745 w_434_604# a_381_614# 0.027639f
C746 a_884_498# p3p2p1g0 0.016011f
C747 g3 p3p2p1p0c0 0.001229f
C748 a_251_466# gnd 0.701773f
C749 a_302_20# a0 0.413834f
C750 w_291_180# a_304_190# 0.019526f
C751 b1 g1 0.281479f
C752 w_758_272# c2 0.003448f
C753 cin vdd 0.057277f
C754 a_397_472# w_450_462# 0.027639f
C755 gnd a3 0.417128f
C756 w_581_n75# a_594_n65# 0.019526f
C757 w_548_n81# a1 0.02809f
C758 w_400_n106# b1 0.015139f
C759 p0 w_693_68# 0.001671f
C760 p1 w_258_n117# 0.013216f
C761 a_239_604# w_226_594# 0.019526f
C762 a_731_417# w_725_411# 0.017071f
C763 vdd a_445_140# 0.41238f
C764 w_367_n112# a_302_n114# 0.015055f
C765 p1g0 p1p0c0 0.011688f
C766 p3p2p1g0 w_877_451# 0.012016f
C767 gnd a_271_280# 0.20619f
C768 w_328_18# vdd 0.001288f
C769 a_380_291# vdd 0.441416f
C770 a_617_278# a_617_318# 0.41238f
C771 w_797_280# vdd 0.001288f
C772 w_834_277# a_847_245# 0.013216f
C773 a_496_251# a_453_311# 0.41238f
C774 p3g2 gnd 0.300358f
C775 p3p2g1 p3p2p1p0c0 0.001238f
C776 p2p1p0c0 a_534_474# 0.060798f
C777 w_658_464# g2 0.005833f
C778 a_534_474# p2g1 9.1e-19
C779 w_854_n201# s2 0.007992f
C780 vdd w_571_625# 0.008451f
C781 a_239_604# a_206_556# 0.003752f
C782 w_347_461# g1 0.01132f
C783 p1 a_594_556# 0.018694f
C784 cin a_797_566# 2.14e-20
C785 g1 a_381_614# 0.059029f
C786 p1 a1 0.008941f
C787 vdd a_617_318# 0.41238f
C788 p0 a_496_232# 0.013746f
C789 vdd gnd 3.54422f
C790 vdd a_795_n247# 0.446951f
C791 a_397_472# vdd 1.32165f
C792 w_367_185# a_380_153# 0.013216f
C793 w_291_180# a_271_142# 0.026794f
C794 a_693_378# w_725_411# 0.013329f
C795 g0 w_611_340# 5.72e-19
C796 c3 a_825_350# 2.29e-19
C797 vdd b2 0.006748f
C798 gnd a_798_n113# 0.206673f
C799 vdd a_269_20# 0.441416f
C800 p3 c3 0.03105f
C801 w_472_604# p3p2g1 0.013216f
C802 w_368_n246# b2 0.01395f
C803 a_738_234# a_771_282# 0.286223f
C804 p1 g1 0.015873f
C805 p0 g2 0.003698f
C806 w_867_n335# p3 0.007896f
C807 a_564_25# gnd 0.20619f
C808 w_504_133# a_445_147# 0.027289f
C809 w_439_134# a_445_140# 0.017071f
C810 gnd s0 0.20619f
C811 p1 w_400_n106# 3.76e-36
C812 cin p2 0.005335f
C813 a_688_664# p3 0.002444f
C814 w_785_n81# vdd 0.030269f
C815 c4 a_825_350# 0.060798f
C816 w_368_n380# b3 0.01395f
C817 w_401_n374# a3 0.028034f
C818 a_324_n46# vdd 0.450999f
C819 vdd pocin 0.440403f
C820 vdd a_302_n114# 0.019283f
C821 g0 c1 0.031415f
C822 a_825_350# w_942_382# 0.027289f
C823 a_883_389# w_877_383# 0.017071f
C824 w_690_n70# vdd 0.008451f
C825 w_834_277# c3 3.18e-20
C826 w_205_450# gnd 2.22e-19
C827 w_473_301# p1g0 0.004305f
C828 p3g2 a_315_567# 0.060798f
C829 c1 a_597_73# 2.15e-19
C830 w_785_n81# a_798_n113# 0.013216f
C831 p3p2g1 a_381_614# 0.060798f
C832 gnd a_239_604# 0.248155f
C833 c3 a_873_n248# 4.29e-20
C834 a_797_547# p3 0.013746f
C835 g3 w_693_n346# 0.013222f
C836 w_328_18# a0 0.007896f
C837 w_658_464# vdd 0.008451f
C838 p2 gnd 1.81974f
C839 a_731_457# a_731_417# 0.41238f
C840 p2 a_795_n247# 0.060798f
C841 a_327_429# g2 0.002808f
C842 a_518_635# w_571_625# 0.027639f
C843 g0 w_604_625# 0.026794f
C844 p2g1 a_610_414# 0.019171f
C845 p0 w_258_174# 0.028034f
C846 p1 g3 0.028063f
C847 p1 a_440_393# 0.013746f
C848 w_401_n374# vdd 0.028764f
C849 p0 a_610_395# 0.019134f
C850 a_594_n65# b1 0.7623f
C851 w_693_n346# a_673_n378# 0.026907f
C852 vdd a_315_567# 0.464809f
C853 a_518_635# gnd 0.042086f
C854 w_367_323# a_304_328# 0.026907f
C855 g2 a2 0.012963f
C856 w_506_301# vdd 0.008451f
C857 p2 a_397_472# 0.002835f
C858 a_847_245# c3 0.006337f
C859 w_581_n75# vdd 2.04e-19
C860 cin p2p1p0c0 0.006726f
C861 gnd a0 1.47749f
C862 p2 b2 0.6987f
C863 cin p2g1 0.013147f
C864 g0 a_534_474# 1.63e-19
C865 a_610_395# a_610_377# 0.41238f
C866 p1 p1g0 7.17e-19
C867 w_400_323# p1g0 0.013216f
C868 p1 p3p2g1 0.017215f
C869 p0 p3g2 0.00253f
C870 p1 c2 0.003604f
C871 cin a_600_239# 8.95e-19
C872 a_688_664# w_675_654# 0.017642f
C873 w_401_604# a_381_614# 0.027639f
C874 a_564_n389# b3 0.00288f
C875 w_434_604# g1 0.026794f
C876 w_795_n349# vdd 0.008639f
C877 w_834_277# a_771_282# 0.027261f
C878 w_439_134# pocin 1.21e-19
C879 a_886_n382# c3 0.002154f
C880 c2 a_816_233# 3.8e-19
C881 w_611_272# p1p0c0 0.057514f
C882 a_424_535# gnd 0.416913f
C883 a_424_554# a_381_614# 0.41238f
C884 g3 p3p2p1g0 0.001198f
C885 a1 g1 0.115698f
C886 a_883_464# a_883_429# 0.41238f
C887 w_725_266# c2 0.003448f
C888 a_397_472# w_417_462# 0.027639f
C889 p0 vdd 0.809918f
C890 a_693_378# w_790_410# 0.027289f
C891 w_440_301# vdd 0.008451f
C892 gnd a_597_n341# 0.701814f
C893 s2 a_873_n248# 0.20619f
C894 w_400_n106# a1 0.028034f
C895 w_367_n112# b1 0.01395f
C896 a_251_466# a_327_429# 0.060798f
C897 a_325_n314# gnd 0.206673f
C898 p0 w_660_68# 0.004686f
C899 a_731_417# w_725_444# 0.008113f
C900 a_883_464# p3p2p1p0c0 0.005542f
C901 p2p1p0c0 gnd 0.207724f
C902 vdd a_445_147# 0.001532f
C903 w_328_n116# a_302_n114# 0.007992f
C904 p2g1 gnd 0.215208f
C905 p3p2g1 w_877_451# 0.037044f
C906 p1g0 a_453_311# 0.010005f
C907 w_291_17# vdd 0.008507f
C908 w_758_272# vdd 6.13e-19
C909 a_847_245# a_771_282# 0.060798f
C910 a_617_278# p1p0c0 0.019123f
C911 p3g2 p3p2p1p0c0 0.001239f
C912 p3p2g1 p3p2p1g0 0.0533f
C913 a_397_472# w_384_462# 0.017642f
C914 gnd a_564_n251# 0.20619f
C915 a_731_457# a_731_492# 0.41238f
C916 p1 s1 0.413834f
C917 p2p1g0 a_534_474# 0.043704f
C918 a_600_239# gnd 0.829424f
C919 w_857_n67# c1 0.027735f
C920 w_620_464# g2 0.00583f
C921 a_397_472# p2g1 0.009943f
C922 gnd a_673_36# 0.248155f
C923 a_808_n381# vdd 0.439903f
C924 a_883_429# vdd 5.02e-19
C925 w_815_n209# s2 0.015055f
C926 vdd w_538_625# 0.008451f
C927 w_314_461# g1 0.01132f
C928 w_347_461# g2 0.005799f
C929 a_239_604# a_315_567# 0.060798f
C930 p3 w_726_513# 4.5e-19
C931 vdd p1p0c0 0.439883f
C932 p1 a_594_n65# 0.004757f
C933 p0 a_564_25# 0.003966f
C934 cin a_738_234# 0.024367f
C935 vdd p3p2p1p0c0 0.460861f
C936 p1 a_496_232# 0.013746f
C937 a_325_n180# a_329_n171# 0.14502f
C938 b2 a_564_n251# 0.002958f
C939 a_304_190# vdd 0.017997f
C940 p3 a_206_556# 0.069923f
C941 w_584_n213# a_564_n251# 0.026794f
C942 a_327_429# vdd 0.441435f
C943 vdd w_505_625# 0.008451f
C944 a_302_20# a_328_97# 0.20619f
C945 w_258_174# a_271_142# 0.013216f
C946 g0 w_544_301# 0.00229f
C947 vdd a2 0.198592f
C948 gnd a_561_n113# 0.20619f
C949 p1 w_554_464# 0.041309f
C950 p3p2p1p0c0 w_878_485# 0.018136f
C951 w_291_n117# vdd 0.008507f
C952 vdd a_324_88# 0.45515f
C953 p2 a_440_412# 0.011867f
C954 w_867_n335# c3 0.027759f
C955 w_551_n219# vdd 0.024509f
C956 w_329_n250# b2 0.027716f
C957 w_368_n246# a2 0.028748f
C958 p1 g2 0.006367f
C959 w_828_n343# p3 0.028748f
C960 w_439_167# a_445_140# 0.008113f
C961 w_439_134# a_445_147# 0.013329f
C962 gnd a_738_234# 0.206673f
C963 a_496_251# a_496_232# 0.41238f
C964 a_876_n114# s1 0.20619f
C965 g2 w_521_464# 0.00583f
C966 p0 p2 0.021182f
C967 cin p3 0.00353f
C968 c3 c1 2.14e-19
C969 w_472_604# vdd 0.008451f
C970 g3 g1 0.023266f
C971 p2p1p0c0 w_658_464# 0.013216f
C972 w_676_271# g1 0.002127f
C973 w_329_n384# b3 0.027716f
C974 w_611_305# a_617_318# 0.009864f
C975 w_368_n380# a3 0.028748f
C976 cin g0 0.023739f
C977 b1 vdd 0.019028f
C978 vdd a_271_142# 0.439904f
C979 a_325_n314# w_401_n374# 0.013216f
C980 p2 a_610_377# 0.013746f
C981 a_693_378# g2 1.39e-20
C982 g0 a_445_140# 0.016231f
C983 p0 a0 0.007613f
C984 a_883_429# a_883_389# 0.41238f
C985 a_883_389# w_877_416# 0.008113f
C986 a_825_350# w_877_383# 0.013329f
C987 p0 w_551_57# 0.00465f
C988 g1 p1g0 0.038781f
C989 g0 a_380_291# 0.008577f
C990 c3 a_771_282# 0.007917f
C991 p3 s3 0.413834f
C992 p3g2 a_381_614# 0.011947f
C993 c2 g1 0.014621f
C994 a_883_389# p3p2p1p0c0 0.016619f
C995 a_825_350# gnd 1.36074f
C996 p2 w_538_625# 0.026794f
C997 c3 s2 0.015855f
C998 w_620_464# vdd 0.008451f
C999 p3 gnd 1.77527f
C1000 a_518_635# w_538_625# 0.027639f
C1001 p1 a_610_395# 0.013746f
C1002 w_845_654# p3p2p1p0c0 0.013216f
C1003 a_594_n65# a1 0.001371f
C1004 w_347_461# vdd 0.008451f
C1005 g0 gnd 0.2831f
C1006 w_291_318# a_304_328# 0.019526f
C1007 vdd a_381_614# 1.32165f
C1008 w_473_301# vdd 0.008451f
C1009 w_548_n81# vdd 0.0086f
C1010 c4 w_942_382# 0.013216f
C1011 cin p2p1g0 0.070233f
C1012 p0 p2p1p0c0 0.00185f
C1013 gnd a_597_73# 0.248155f
C1014 p2 a2 0.49284f
C1015 p0 p2g1 0.007444f
C1016 g0 a_397_472# 0.059421f
C1017 a_518_635# w_505_625# 0.017642f
C1018 p1 a_271_280# 0.060798f
C1019 a_797_604# a_797_585# 0.41238f
C1020 p1 p3g2 0.057343f
C1021 g3 a_673_n378# 0.060798f
C1022 a_884_498# a_883_464# 0.41238f
C1023 p0 a_673_36# 0.003088f
C1024 p1 w_741_654# 0.026794f
C1025 w_657_n70# a_670_n102# 0.013216f
C1026 a_564_n389# a3 0.060856f
C1027 w_368_604# a_381_614# 0.017642f
C1028 w_335_599# a_315_567# 0.026907f
C1029 w_581_n75# a_561_n113# 0.026794f
C1030 w_693_n346# vdd 0.008611f
C1031 w_439_167# pocin 0.036563f
C1032 a_304_328# a_271_280# 0.003752f
C1033 a_886_n382# 0 0.016528f $  
C1034 s3 0 0.473154f $  
C1035 a_808_n381# 0 0.526842f $  
C1036 a_564_n389# 0 0.477455f $  
C1037 a_673_n378# 0 0.382299f $  
C1038 a_329_n305# 0 0.016528f $  
C1039 a_325_n314# 0 0.526842f $  
C1040 b3 0 6.62907f $  
C1041 a3 0 2.45012f $  
C1042 a_597_n341# 0 0.771781f $  
C1043 a_873_n248# 0 0.016528f $  
C1044 s2 0 0.462937f $  
C1045 a_795_n247# 0 0.526842f $  
C1046 a_564_n251# 0 0.477455f $  
C1047 a_329_n171# 0 0.016528f $  
C1048 a_325_n180# 0 0.526842f $  
C1049 b2 0 6.55321f $  
C1050 a2 0 2.34823f $  
C1051 a_876_n114# 0 0.016528f $  
C1052 s1 0 0.462937f $  
C1053 a_798_n113# 0 0.526842f $  
C1054 a_561_n113# 0 0.477455f $  
C1055 a_670_n102# 0 0.382299f $  
C1056 a_328_n37# 0 0.016528f $  
C1057 a_302_n114# 0 0.662497f $  
C1058 a_269_n114# 0 0.382299f $  
C1059 a_324_n46# 0 0.526842f $  
C1060 b1 0 5.67351f $  
C1061 a1 0 2.3497f $  
C1062 a_594_n65# 0 0.771781f $  
C1063 a_564_25# 0 0.477455f $  
C1064 a_673_36# 0 0.382299f $  
C1065 a_328_97# 0 0.016528f $  
C1066 a_302_20# 0 0.662497f $  
C1067 a_269_20# 0 0.382299f $  
C1068 a_324_88# 0 0.526842f $  
C1069 b0 0 6.55052f $  
C1070 a0 0 2.47333f $  
C1071 a_597_73# 0 0.804448f $  
C1072 c1 0 2.23371f $  
C1073 a_445_140# 0 0.179875f $  
C1074 a_445_147# 0 1.02677f $  
C1075 a_816_233# 0 0.016528f $  
C1076 pocin 0 0.599293f $  
C1077 a_271_142# 0 0.477455f $  
C1078 a_380_153# 0 0.382299f $  
C1079 a_496_232# 0 0.040245f $  
C1080 s0 0 0.145867f $  
C1081 a_738_234# 0 0.526842f $  
C1082 a_304_190# 0 0.771781f $  
C1083 a_496_251# 0 0.040245f $  
C1084 c2 0 2.27948f $  
C1085 a_617_278# 0 0.206277f $  
C1086 a_600_239# 0 1.28245f $  
C1087 a_847_245# 0 0.382299f $  
C1088 a_771_282# 0 0.662497f $  
C1089 a_617_318# 0 0.150155f $  
C1090 p1p0c0 0 0.596493f $  
C1091 a_453_311# 0 1.70512f $  
C1092 p1g0 0 1.48359f $  
C1093 a_271_280# 0 0.477455f $  
C1094 c4 0 0.147767f $  
C1095 a_380_291# 0 0.382299f $  
C1096 a_610_377# 0 0.036687f $  
C1097 a_304_328# 0 0.771914f $  
C1098 a_440_393# 0 0.040245f $  
C1099 a_610_395# 0 0.040245f $  
C1100 a_883_389# 0 0.206277f $  
C1101 a_825_350# 0 1.81542f $  
C1102 c3 0 2.59712f $  
C1103 a_610_414# 0 0.040245f $  
C1104 a_440_412# 0 0.040245f $  
C1105 a_731_417# 0 0.206277f $  
C1106 a_883_429# 0 0.150155f $  
C1107 a_693_378# 0 1.54889f $  
C1108 a_731_457# 0 0.150155f $  
C1109 a_883_464# 0 0.148414f $  
C1110 p2p1p0c0 0 1.71192f $  
C1111 p2p1g0 0 1.59696f $  
C1112 p2g1 0 0.842448f $  
C1113 a_218_418# 0 0.477455f $  
C1114 a_534_474# 0 2.13082f $  
C1115 a_397_472# 0 1.70506f $  
C1116 a_327_429# 0 0.382299f $  
C1117 a_731_492# 0 0.148414f $  
C1118 a_884_498# 0 0.144831f $  
C1119 g3 0 6.00295f $  
C1120 a_251_466# 0 0.770807f $  
C1121 a_424_535# 0 0.040245f $  
C1122 a_594_537# 0 0.040245f $  
C1123 a_797_547# 0 0.040245f $  
C1124 a_594_556# 0 0.040245f $  
C1125 a_424_554# 0 0.040245f $  
C1126 a_797_566# 0 0.040245f $  
C1127 a_594_575# 0 0.040245f $  
C1128 a_797_585# 0 0.040245f $  
C1129 a_797_604# 0 0.040245f $  
C1130 gnd 0 32.550102f $  
C1131 p3p2p1p0c0 0 4.09846f $  
C1132 p3p2p1g0 0 6.27811f $  
C1133 p3p2g1 0 4.70971f $  
C1134 p3g2 0 5.74969f $  
C1135 vdd 0 38.531303f $  
C1136 a_206_556# 0 0.477455f $  
C1137 a_315_567# 0 0.382299f $  
C1138 a_381_614# 0 1.70511f $  
C1139 g1 0 21.4853f $  
C1140 g2 0 19.795301f $  
C1141 a_239_604# 0 0.804448f $  
C1142 a_518_635# 0 2.1423f $  
C1143 g0 0 15.508599f $  
C1144 a_688_664# 0 2.57948f $  
C1145 cin 0 4.54177f $  
C1146 p0 0 7.20932f $  
C1147 p1 0 13.8549f $  
C1148 p2 0 13.4502f $  
C1149 p3 0 14.974599f $  
C1150 w_867_n335# 0 1.25349f $  
C1151 w_828_n343# 0 1.34991f $  
C1152 w_795_n349# 0 1.34991f $  
C1153 w_693_n346# 0 1.34991f $  
C1154 w_660_n346# 0 1.34991f $  
C1155 w_584_n351# 0 1.34991f $  
C1156 w_551_n357# 0 1.34991f $  
C1157 w_401_n374# 0 1.34991f $  
C1158 w_368_n380# 0 1.34991f $  
C1159 w_329_n384# 0 1.25349f $  
C1160 w_854_n201# 0 1.25349f $  
C1161 w_815_n209# 0 1.34991f $  
C1162 w_782_n215# 0 1.34991f $  
C1163 w_584_n213# 0 1.34991f $  
C1164 w_551_n219# 0 1.34991f $  
C1165 w_401_n240# 0 1.34991f $  
C1166 w_368_n246# 0 1.34991f $  
C1167 w_329_n250# 0 1.25349f $  
C1168 w_857_n67# 0 1.25349f $  
C1169 w_818_n75# 0 1.34991f $  
C1170 w_785_n81# 0 1.34991f $  
C1171 w_690_n70# 0 1.34991f $  
C1172 w_657_n70# 0 1.34991f $  
C1173 w_581_n75# 0 1.34991f $  
C1174 w_548_n81# 0 1.34991f $  
C1175 w_400_n106# 0 1.34991f $  
C1176 w_367_n112# 0 1.34991f $  
C1177 w_328_n116# 0 1.25349f $  
C1178 w_291_n117# 0 1.34991f $  
C1179 w_258_n117# 0 1.34991f $  
C1180 w_693_68# 0 1.34991f $  
C1181 w_660_68# 0 1.34991f $  
C1182 w_584_63# 0 1.34991f $  
C1183 w_551_57# 0 1.34991f $  
C1184 w_400_28# 0 1.34991f $  
C1185 w_367_22# 0 1.34991f $  
C1186 w_328_18# 0 1.25349f $  
C1187 w_291_17# 0 1.34991f $  
C1188 w_258_17# 0 1.34991f $  
C1189 w_504_133# 0 1.34991f $  
C1190 w_439_134# 0 1.34991f $  
C1191 w_439_167# 0 1.34991f $  
C1192 w_400_185# 0 1.34991f $  
C1193 w_367_185# 0 1.34991f $  
C1194 w_291_180# 0 1.34991f $  
C1195 w_258_174# 0 1.34991f $  
C1196 w_867_277# 0 1.34991f $  
C1197 w_834_277# 0 1.34991f $  
C1198 w_797_280# 0 1.25349f $  
C1199 w_758_272# 0 1.34991f $  
C1200 w_725_266# 0 1.34991f $  
C1201 w_676_271# 0 1.34991f $  
C1202 w_611_272# 0 1.34991f $  
C1203 w_611_305# 0 1.34991f $  
C1204 w_611_340# 0 1.34991f $  
C1205 w_544_301# 0 1.34991f $  
C1206 w_506_301# 0 1.34991f $  
C1207 w_473_301# 0 1.34991f $  
C1208 w_440_301# 0 1.34991f $  
C1209 w_400_323# 0 1.34991f $  
C1210 w_367_323# 0 1.34991f $  
C1211 w_291_318# 0 1.34991f $  
C1212 w_258_312# 0 1.34991f $  
C1213 w_942_382# 0 1.34991f $  
C1214 w_877_383# 0 1.34991f $  
C1215 w_877_416# 0 1.34991f $  
C1216 w_877_451# 0 1.34991f $  
C1217 w_790_410# 0 1.34991f $  
C1218 w_725_411# 0 1.34991f $  
C1219 w_725_444# 0 1.34991f $  
C1220 w_878_485# 0 1.34991f $  
C1221 w_725_479# 0 1.34991f $  
C1222 w_879_518# 0 1.34991f $  
C1223 w_726_513# 0 1.34991f $  
C1224 w_658_464# 0 1.34991f $  
C1225 w_620_464# 0 1.34991f $  
C1226 w_587_464# 0 1.34991f $  
C1227 w_554_464# 0 1.34991f $  
C1228 w_521_464# 0 1.34991f $  
C1229 w_488_462# 0 1.34991f $  
C1230 w_450_462# 0 1.34991f $  
C1231 w_417_462# 0 1.34991f $  
C1232 w_384_462# 0 1.34991f $  
C1233 w_347_461# 0 1.34991f $  
C1234 w_314_461# 0 1.34991f $  
C1235 w_238_456# 0 1.34991f $  
C1236 w_205_450# 0 1.34991f $  
C1237 w_845_654# 0 1.34991f $  
C1238 w_807_654# 0 1.34991f $  
C1239 w_774_654# 0 1.34991f $  
C1240 w_741_654# 0 1.34991f $  
C1241 w_708_654# 0 1.34991f $  
C1242 w_675_654# 0 1.34991f $  
C1243 w_642_625# 0 1.34991f $  
C1244 w_604_625# 0 1.34991f $  
C1245 w_571_625# 0 1.34991f $  
C1246 w_538_625# 0 1.34991f $  
C1247 w_505_625# 0 1.34991f $  
C1248 w_472_604# 0 1.34991f $  
C1249 w_434_604# 0 1.34991f $  
C1250 w_401_604# 0 1.34991f $  
C1251 w_368_604# 0 1.34991f $  
C1252 w_335_599# 0 1.34991f $  
C1253 w_302_599# 0 1.34991f $  
C1254 w_226_594# 0 1.34991f $  
C1255 w_193_588# 0 1.34991f $  










 

* * RISING AND FALLING DELAY MEASUREMENT
* * * Measure the delay for the final carry-out signal (C4)
.measure tran delay_C4_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(c4) VAL=0.9 FALL=1
.measure tran delay_C4_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(c4) VAL=0.9 RISE=1

* * Measure the delay for each sum signal
.measure tran delay_S0_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s0) VAL=0.9 FALL=1
.measure tran delay_S0_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s0) VAL=0.9 RISE=1
.measure tran delay_S1_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s1) VAL=0.9 FALL=1
.measure tran delay_S1_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s1) VAL=0.9 RISE=1
.measure tran delay_S2_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s2) VAL=0.9 FALL=1
.measure tran delay_S2_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s2) VAL=0.9 RISE=1
.measure tran delay_S3_fall TRIG V(a0) VAL=0.9 FALL=1 TARG V(s3) VAL=0.9 FALL=1
.measure tran delay_S3_rise TRIG V(a0) VAL=0.9 RISE=1 TARG V(s3) VAL=0.9 RISE=1



.control
  set hcopypscolor = 1             
  set color0 = white               
  set color1 = black               
  set color2 = red                 
  set color3 = blue                
  set color4 = coral               
  set color5 = brown    
  set color6 = cyan
  set color7 = chocolate   
  set color8 = chocolate
  set color9 = blueviolet
  set color10 = cadetblue        
  * for testing        
  * tran 1n 160n
  * for delay  
  tran 0.01n 40n 
   plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+g0 20+g1 22+g2 24+g3   
  plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+p0 20+p1 22+p2 24+p3                      
  * plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+s0 20+s1 22+s2 24+s3                      
    plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+c4 20+s0 22+s1 24+s2 26+s3   
    plot pocin 2+g0 4+c1
    * plot g3 2+p3g2 4+p3p2g1 6+p3p2p1g0 8+p3p2p1p0c0 10+c4 
    plot c1 2+p1 4+s1
  plot s0 2+s1 4+s2 6+s3    
        
.endc