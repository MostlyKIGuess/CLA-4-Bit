* OR Testing Code
* TSMC 180nm Technology Parameters
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* Test Signals
Vclk b gnd PULSE(0 'SUPPLY' 0 0.001n 0.01n 10n 20n)
Vd c gnd PULSE(0 'SUPPLY' 0n 0.001n 0.01n 35n 70n)

* SPICE3 file created from or.ext - technology: scmos
.option scale=0.09u

M1000 ybar b gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 ybar c gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 ybar c a_n75_7# w_n81_1# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1003 y ybar vdd w_n16_0# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 vdd b a_n75_7# w_n81_34# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1005 y ybar gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
C0 w_n81_34# vdd 1.41f
C1 gnd ybar 0.808f
C2 w_n81_1# a_n75_7# 2.444f
C3 w_n16_0# vdd 1.128f
C4 c w_n81_1# 2.312f
C5 ybar w_n16_0# 1.014f
C6 w_n81_34# a_n75_7# 1.128f
C7 w_n16_0# y 1.88f
C8 w_n81_34# b 1.482f
C9 w_n81_1# ybar 1.88f
C10 gnd 0 11.561999f 
C11 y 0 4.324f 
C12 c 0 8.299999f 
C13 a_n75_7# 0 4.888f 
C14 b 0 24.082f 
C15 ybar 0 19.995f 
C16 vdd 0 13.536f 

.control
  set hcopypscolor = 1
  set color0 = white
  set color1 = black
  set color2 = red
  set color3 = blue
  set color4 = brown
  set color5 = magenta
  set color6 = cyan
  set color7 = green
  tran 1n 200n
    plot c 2+b 4+y
.endc


