magic
tech scmos
timestamp 1731317385
<< nwell >>
rect 193 588 217 644
rect 226 594 250 650
rect 302 599 326 655
rect 335 599 359 655
rect 368 604 392 660
rect 401 604 425 660
rect 434 604 458 660
rect 472 604 496 660
rect 505 625 529 681
rect 538 625 562 681
rect 571 625 595 681
rect 604 625 628 681
rect 642 625 666 681
rect 675 654 699 710
rect 708 654 732 710
rect 741 654 765 710
rect 774 654 798 710
rect 807 654 831 710
rect 845 654 869 710
rect 205 450 229 506
rect 238 456 262 512
rect 314 461 338 517
rect 347 461 371 517
rect 384 462 408 518
rect 417 462 441 518
rect 450 462 474 518
rect 488 462 512 518
rect 521 464 545 520
rect 554 464 578 520
rect 587 464 611 520
rect 620 464 644 520
rect 658 464 682 520
rect 726 513 782 537
rect 879 518 935 542
rect 725 479 781 503
rect 878 485 934 509
rect 725 444 781 468
rect 725 411 781 435
rect 790 410 814 466
rect 877 451 933 475
rect 877 416 933 440
rect 877 383 933 407
rect 942 382 966 438
rect 258 312 282 368
rect 291 318 315 374
rect 367 323 391 379
rect 400 323 424 379
rect 440 301 464 357
rect 473 301 497 357
rect 506 301 530 357
rect 544 301 568 357
rect 611 340 667 364
rect 611 305 667 329
rect 611 272 667 296
rect 676 271 700 327
rect 725 266 749 322
rect 758 272 782 328
rect 797 280 821 332
rect 834 277 858 333
rect 867 277 891 333
rect 258 174 282 230
rect 291 180 315 236
rect 367 185 391 241
rect 400 185 424 241
rect 439 167 495 191
rect 439 134 495 158
rect 504 133 528 189
rect 258 17 282 73
rect 291 17 315 73
rect 328 18 352 70
rect 367 22 391 78
rect 400 28 424 84
rect 569 57 593 113
rect 602 63 626 119
rect 688 103 712 159
rect 721 109 745 165
rect 760 117 784 169
rect 797 114 821 170
rect 830 114 854 170
rect 258 -117 282 -61
rect 291 -117 315 -61
rect 328 -116 352 -64
rect 367 -112 391 -56
rect 400 -106 424 -50
rect 566 -81 590 -25
rect 599 -75 623 -19
rect 687 -43 711 13
rect 720 -37 744 19
rect 759 -29 783 23
rect 796 -32 820 24
rect 829 -32 853 24
rect 259 -251 283 -195
rect 292 -251 316 -195
rect 329 -250 353 -198
rect 368 -246 392 -190
rect 401 -240 425 -184
rect 569 -219 593 -163
rect 602 -213 626 -157
rect 692 -177 716 -121
rect 725 -171 749 -115
rect 764 -163 788 -111
rect 801 -166 825 -110
rect 834 -166 858 -110
rect 259 -385 283 -329
rect 292 -385 316 -329
rect 329 -384 353 -332
rect 368 -380 392 -324
rect 401 -374 425 -318
rect 569 -357 593 -301
rect 602 -351 626 -295
<< ntransistor >>
rect 252 667 272 669
rect 797 621 837 623
rect 856 622 858 642
rect 252 581 272 583
rect 204 556 206 576
rect 313 567 315 587
rect 346 567 348 587
rect 424 571 464 573
rect 483 572 485 592
rect 594 592 634 594
rect 653 593 655 613
rect 797 602 837 604
rect 797 583 837 585
rect 594 573 634 575
rect 797 564 837 566
rect 424 552 464 554
rect 594 554 634 556
rect 797 545 837 547
rect 424 533 464 535
rect 594 535 634 537
rect 264 529 284 531
rect 264 443 284 445
rect 216 418 218 438
rect 325 429 327 449
rect 358 429 360 449
rect 440 429 480 431
rect 499 430 501 450
rect 610 431 650 433
rect 669 432 671 452
rect 440 410 480 412
rect 610 412 650 414
rect 317 391 337 393
rect 440 391 480 393
rect 610 393 650 395
rect 691 378 693 398
rect 712 378 714 398
rect 741 378 743 398
rect 774 378 776 398
rect 801 378 803 398
rect 610 375 650 377
rect 823 350 825 370
rect 843 350 845 370
rect 864 350 866 370
rect 893 350 895 370
rect 926 350 928 370
rect 953 350 955 370
rect 317 305 337 307
rect 269 280 271 300
rect 378 291 380 311
rect 411 291 413 311
rect 496 268 536 270
rect 555 269 557 289
rect 317 253 337 255
rect 496 249 536 251
rect 598 239 600 259
rect 627 239 629 259
rect 660 239 662 259
rect 687 239 689 259
rect 784 258 804 260
rect 736 234 738 254
rect 496 230 536 232
rect 821 233 823 253
rect 845 245 847 265
rect 878 245 880 265
rect 317 167 337 169
rect 269 142 271 162
rect 378 153 380 173
rect 411 153 413 173
rect 628 136 648 138
rect 269 85 271 105
rect 302 85 304 105
rect 326 97 328 117
rect 411 96 413 116
rect 455 101 457 121
rect 488 101 490 121
rect 515 101 517 121
rect 345 90 365 92
rect 747 95 767 97
rect 699 71 701 91
rect 784 70 786 90
rect 808 82 810 102
rect 841 82 843 102
rect 628 50 648 52
rect 580 25 582 45
rect 625 -2 645 0
rect 269 -49 271 -29
rect 302 -49 304 -29
rect 326 -37 328 -17
rect 411 -38 413 -18
rect 345 -44 365 -42
rect 746 -51 766 -49
rect 698 -75 700 -55
rect 783 -76 785 -56
rect 807 -64 809 -44
rect 840 -64 842 -44
rect 625 -88 645 -86
rect 577 -113 579 -93
rect 628 -140 648 -138
rect 270 -183 272 -163
rect 303 -183 305 -163
rect 327 -171 329 -151
rect 412 -172 414 -152
rect 346 -178 366 -176
rect 751 -185 771 -183
rect 703 -209 705 -189
rect 788 -210 790 -190
rect 812 -198 814 -178
rect 845 -198 847 -178
rect 628 -226 648 -224
rect 580 -251 582 -231
rect 628 -278 648 -276
rect 270 -317 272 -297
rect 303 -317 305 -297
rect 327 -305 329 -285
rect 412 -306 414 -286
rect 346 -312 366 -310
rect 628 -364 648 -362
rect 580 -389 582 -369
<< ptransistor >>
rect 204 598 206 638
rect 237 604 239 644
rect 313 609 315 649
rect 346 609 348 649
rect 379 614 381 654
rect 412 614 414 654
rect 445 614 447 654
rect 483 614 485 654
rect 516 635 518 675
rect 549 635 551 675
rect 582 635 584 675
rect 615 635 617 675
rect 653 635 655 675
rect 686 664 688 704
rect 719 664 721 704
rect 752 664 754 704
rect 785 664 787 704
rect 818 664 820 704
rect 856 664 858 704
rect 885 529 925 531
rect 732 524 772 526
rect 216 460 218 500
rect 249 466 251 506
rect 325 471 327 511
rect 358 471 360 511
rect 395 472 397 512
rect 428 472 430 512
rect 461 472 463 512
rect 499 472 501 512
rect 532 474 534 514
rect 565 474 567 514
rect 598 474 600 514
rect 631 474 633 514
rect 669 474 671 514
rect 884 496 924 498
rect 731 490 771 492
rect 883 462 923 464
rect 731 455 771 457
rect 731 422 771 424
rect 801 420 803 460
rect 883 427 923 429
rect 883 394 923 396
rect 953 392 955 432
rect 269 322 271 362
rect 302 328 304 368
rect 378 333 380 373
rect 411 333 413 373
rect 451 311 453 351
rect 484 311 486 351
rect 517 311 519 351
rect 555 311 557 351
rect 617 351 657 353
rect 617 316 657 318
rect 617 283 657 285
rect 687 281 689 321
rect 736 276 738 316
rect 769 282 771 322
rect 808 286 810 326
rect 845 287 847 327
rect 878 287 880 327
rect 269 184 271 224
rect 302 190 304 230
rect 378 195 380 235
rect 411 195 413 235
rect 445 178 485 180
rect 445 145 485 147
rect 515 143 517 183
rect 699 113 701 153
rect 732 119 734 159
rect 771 123 773 163
rect 808 124 810 164
rect 841 124 843 164
rect 269 23 271 63
rect 302 23 304 63
rect 339 24 341 64
rect 378 28 380 68
rect 411 34 413 74
rect 580 67 582 107
rect 613 73 615 113
rect 269 -111 271 -71
rect 302 -111 304 -71
rect 339 -110 341 -70
rect 378 -106 380 -66
rect 411 -100 413 -60
rect 577 -71 579 -31
rect 610 -65 612 -25
rect 698 -33 700 7
rect 731 -27 733 13
rect 770 -23 772 17
rect 807 -22 809 18
rect 840 -22 842 18
rect 270 -245 272 -205
rect 303 -245 305 -205
rect 340 -244 342 -204
rect 379 -240 381 -200
rect 412 -234 414 -194
rect 580 -209 582 -169
rect 613 -203 615 -163
rect 703 -167 705 -127
rect 736 -161 738 -121
rect 775 -157 777 -117
rect 812 -156 814 -116
rect 845 -156 847 -116
rect 270 -379 272 -339
rect 303 -379 305 -339
rect 340 -378 342 -338
rect 379 -374 381 -334
rect 412 -368 414 -328
rect 580 -347 582 -307
rect 613 -341 615 -301
<< ndiffusion >>
rect 252 669 272 670
rect 252 666 272 667
rect 797 623 837 624
rect 855 622 856 642
rect 858 622 859 642
rect 797 620 837 621
rect 252 583 272 584
rect 252 580 272 581
rect 203 556 204 576
rect 206 556 207 576
rect 312 567 313 587
rect 315 567 316 587
rect 345 567 346 587
rect 348 567 349 587
rect 424 573 464 574
rect 482 572 483 592
rect 485 572 486 592
rect 594 594 634 595
rect 652 593 653 613
rect 655 593 656 613
rect 797 604 837 605
rect 797 601 837 602
rect 594 591 634 592
rect 797 585 837 586
rect 797 582 837 583
rect 424 570 464 571
rect 594 575 634 576
rect 594 572 634 573
rect 797 566 837 567
rect 797 563 837 564
rect 424 554 464 555
rect 594 556 634 557
rect 594 553 634 554
rect 424 551 464 552
rect 797 547 837 548
rect 797 544 837 545
rect 264 531 284 532
rect 424 535 464 536
rect 594 537 634 538
rect 594 534 634 535
rect 424 532 464 533
rect 264 528 284 529
rect 264 445 284 446
rect 264 442 284 443
rect 215 418 216 438
rect 218 418 219 438
rect 324 429 325 449
rect 327 429 328 449
rect 357 429 358 449
rect 360 429 361 449
rect 440 431 480 432
rect 498 430 499 450
rect 501 430 502 450
rect 440 428 480 429
rect 610 433 650 434
rect 668 432 669 452
rect 671 432 672 452
rect 610 430 650 431
rect 440 412 480 413
rect 610 414 650 415
rect 610 411 650 412
rect 440 409 480 410
rect 317 393 337 394
rect 317 390 337 391
rect 440 393 480 394
rect 610 395 650 396
rect 610 392 650 393
rect 440 390 480 391
rect 690 378 691 398
rect 693 378 694 398
rect 711 378 712 398
rect 714 378 715 398
rect 740 378 741 398
rect 743 378 744 398
rect 773 378 774 398
rect 776 378 777 398
rect 800 378 801 398
rect 803 378 804 398
rect 610 377 650 378
rect 610 374 650 375
rect 822 350 823 370
rect 825 350 826 370
rect 842 350 843 370
rect 845 350 846 370
rect 863 350 864 370
rect 866 350 867 370
rect 892 350 893 370
rect 895 350 896 370
rect 925 350 926 370
rect 928 350 929 370
rect 952 350 953 370
rect 955 350 956 370
rect 317 307 337 308
rect 317 304 337 305
rect 268 280 269 300
rect 271 280 272 300
rect 377 291 378 311
rect 380 291 381 311
rect 410 291 411 311
rect 413 291 414 311
rect 496 270 536 271
rect 554 269 555 289
rect 557 269 558 289
rect 496 267 536 268
rect 317 255 337 256
rect 317 252 337 253
rect 496 251 536 252
rect 496 248 536 249
rect 597 239 598 259
rect 600 239 601 259
rect 626 239 627 259
rect 629 239 630 259
rect 659 239 660 259
rect 662 239 663 259
rect 686 239 687 259
rect 689 239 690 259
rect 784 260 804 261
rect 784 257 804 258
rect 735 234 736 254
rect 738 234 739 254
rect 496 232 536 233
rect 820 233 821 253
rect 823 233 824 253
rect 844 245 845 265
rect 847 245 848 265
rect 877 245 878 265
rect 880 245 881 265
rect 496 229 536 230
rect 317 169 337 170
rect 317 166 337 167
rect 268 142 269 162
rect 271 142 272 162
rect 377 153 378 173
rect 380 153 381 173
rect 410 153 411 173
rect 413 153 414 173
rect 628 138 648 139
rect 628 135 648 136
rect 268 85 269 105
rect 271 85 272 105
rect 301 85 302 105
rect 304 85 305 105
rect 325 97 326 117
rect 328 97 329 117
rect 410 96 411 116
rect 413 96 414 116
rect 454 101 455 121
rect 457 101 458 121
rect 487 101 488 121
rect 490 101 491 121
rect 514 101 515 121
rect 517 101 518 121
rect 345 92 365 93
rect 345 89 365 90
rect 747 97 767 98
rect 747 94 767 95
rect 698 71 699 91
rect 701 71 702 91
rect 783 70 784 90
rect 786 70 787 90
rect 807 82 808 102
rect 810 82 811 102
rect 840 82 841 102
rect 843 82 844 102
rect 628 52 648 53
rect 628 49 648 50
rect 579 25 580 45
rect 582 25 583 45
rect 625 0 645 1
rect 625 -3 645 -2
rect 268 -49 269 -29
rect 271 -49 272 -29
rect 301 -49 302 -29
rect 304 -49 305 -29
rect 325 -37 326 -17
rect 328 -37 329 -17
rect 410 -38 411 -18
rect 413 -38 414 -18
rect 345 -42 365 -41
rect 345 -45 365 -44
rect 746 -49 766 -48
rect 746 -52 766 -51
rect 697 -75 698 -55
rect 700 -75 701 -55
rect 782 -76 783 -56
rect 785 -76 786 -56
rect 806 -64 807 -44
rect 809 -64 810 -44
rect 839 -64 840 -44
rect 842 -64 843 -44
rect 625 -86 645 -85
rect 625 -89 645 -88
rect 576 -113 577 -93
rect 579 -113 580 -93
rect 628 -138 648 -137
rect 628 -141 648 -140
rect 269 -183 270 -163
rect 272 -183 273 -163
rect 302 -183 303 -163
rect 305 -183 306 -163
rect 326 -171 327 -151
rect 329 -171 330 -151
rect 411 -172 412 -152
rect 414 -172 415 -152
rect 346 -176 366 -175
rect 346 -179 366 -178
rect 751 -183 771 -182
rect 751 -186 771 -185
rect 702 -209 703 -189
rect 705 -209 706 -189
rect 787 -210 788 -190
rect 790 -210 791 -190
rect 811 -198 812 -178
rect 814 -198 815 -178
rect 844 -198 845 -178
rect 847 -198 848 -178
rect 628 -224 648 -223
rect 628 -227 648 -226
rect 579 -251 580 -231
rect 582 -251 583 -231
rect 628 -276 648 -275
rect 628 -279 648 -278
rect 269 -317 270 -297
rect 272 -317 273 -297
rect 302 -317 303 -297
rect 305 -317 306 -297
rect 326 -305 327 -285
rect 329 -305 330 -285
rect 411 -306 412 -286
rect 414 -306 415 -286
rect 346 -310 366 -309
rect 346 -313 366 -312
rect 628 -362 648 -361
rect 628 -365 648 -364
rect 579 -389 580 -369
rect 582 -389 583 -369
<< pdiffusion >>
rect 203 598 204 638
rect 206 598 207 638
rect 236 604 237 644
rect 239 604 240 644
rect 312 609 313 649
rect 315 609 316 649
rect 345 609 346 649
rect 348 609 349 649
rect 378 614 379 654
rect 381 614 382 654
rect 411 614 412 654
rect 414 614 415 654
rect 444 614 445 654
rect 447 614 448 654
rect 482 614 483 654
rect 485 614 486 654
rect 515 635 516 675
rect 518 635 519 675
rect 548 635 549 675
rect 551 635 552 675
rect 581 635 582 675
rect 584 635 585 675
rect 614 635 615 675
rect 617 635 618 675
rect 652 635 653 675
rect 655 635 656 675
rect 685 664 686 704
rect 688 664 689 704
rect 718 664 719 704
rect 721 664 722 704
rect 751 664 752 704
rect 754 664 755 704
rect 784 664 785 704
rect 787 664 788 704
rect 817 664 818 704
rect 820 664 821 704
rect 855 664 856 704
rect 858 664 859 704
rect 885 531 925 532
rect 885 528 925 529
rect 732 526 772 527
rect 732 523 772 524
rect 215 460 216 500
rect 218 460 219 500
rect 248 466 249 506
rect 251 466 252 506
rect 324 471 325 511
rect 327 471 328 511
rect 357 471 358 511
rect 360 471 361 511
rect 394 472 395 512
rect 397 472 398 512
rect 427 472 428 512
rect 430 472 431 512
rect 460 472 461 512
rect 463 472 464 512
rect 498 472 499 512
rect 501 472 502 512
rect 531 474 532 514
rect 534 474 535 514
rect 564 474 565 514
rect 567 474 568 514
rect 597 474 598 514
rect 600 474 601 514
rect 630 474 631 514
rect 633 474 634 514
rect 668 474 669 514
rect 671 474 672 514
rect 884 498 924 499
rect 884 495 924 496
rect 731 492 771 493
rect 731 489 771 490
rect 883 464 923 465
rect 883 461 923 462
rect 731 457 771 458
rect 731 454 771 455
rect 731 424 771 425
rect 731 421 771 422
rect 800 420 801 460
rect 803 420 804 460
rect 883 429 923 430
rect 883 426 923 427
rect 883 396 923 397
rect 883 393 923 394
rect 952 392 953 432
rect 955 392 956 432
rect 268 322 269 362
rect 271 322 272 362
rect 301 328 302 368
rect 304 328 305 368
rect 377 333 378 373
rect 380 333 381 373
rect 410 333 411 373
rect 413 333 414 373
rect 450 311 451 351
rect 453 311 454 351
rect 483 311 484 351
rect 486 311 487 351
rect 516 311 517 351
rect 519 311 520 351
rect 554 311 555 351
rect 557 311 558 351
rect 617 353 657 354
rect 617 350 657 351
rect 617 318 657 319
rect 617 315 657 316
rect 617 285 657 286
rect 617 282 657 283
rect 686 281 687 321
rect 689 281 690 321
rect 735 276 736 316
rect 738 276 739 316
rect 768 282 769 322
rect 771 282 772 322
rect 807 286 808 326
rect 810 286 811 326
rect 844 287 845 327
rect 847 287 848 327
rect 877 287 878 327
rect 880 287 881 327
rect 268 184 269 224
rect 271 184 272 224
rect 301 190 302 230
rect 304 190 305 230
rect 377 195 378 235
rect 380 195 381 235
rect 410 195 411 235
rect 413 195 414 235
rect 445 180 485 181
rect 445 177 485 178
rect 445 147 485 148
rect 445 144 485 145
rect 514 143 515 183
rect 517 143 518 183
rect 698 113 699 153
rect 701 113 702 153
rect 731 119 732 159
rect 734 119 735 159
rect 770 123 771 163
rect 773 123 774 163
rect 807 124 808 164
rect 810 124 811 164
rect 840 124 841 164
rect 843 124 844 164
rect 268 23 269 63
rect 271 23 272 63
rect 301 23 302 63
rect 304 23 305 63
rect 338 24 339 64
rect 341 24 342 64
rect 377 28 378 68
rect 380 28 381 68
rect 410 34 411 74
rect 413 34 414 74
rect 579 67 580 107
rect 582 67 583 107
rect 612 73 613 113
rect 615 73 616 113
rect 268 -111 269 -71
rect 271 -111 272 -71
rect 301 -111 302 -71
rect 304 -111 305 -71
rect 338 -110 339 -70
rect 341 -110 342 -70
rect 377 -106 378 -66
rect 380 -106 381 -66
rect 410 -100 411 -60
rect 413 -100 414 -60
rect 576 -71 577 -31
rect 579 -71 580 -31
rect 609 -65 610 -25
rect 612 -65 613 -25
rect 697 -33 698 7
rect 700 -33 701 7
rect 730 -27 731 13
rect 733 -27 734 13
rect 769 -23 770 17
rect 772 -23 773 17
rect 806 -22 807 18
rect 809 -22 810 18
rect 839 -22 840 18
rect 842 -22 843 18
rect 269 -245 270 -205
rect 272 -245 273 -205
rect 302 -245 303 -205
rect 305 -245 306 -205
rect 339 -244 340 -204
rect 342 -244 343 -204
rect 378 -240 379 -200
rect 381 -240 382 -200
rect 411 -234 412 -194
rect 414 -234 415 -194
rect 579 -209 580 -169
rect 582 -209 583 -169
rect 612 -203 613 -163
rect 615 -203 616 -163
rect 702 -167 703 -127
rect 705 -167 706 -127
rect 735 -161 736 -121
rect 738 -161 739 -121
rect 774 -157 775 -117
rect 777 -157 778 -117
rect 811 -156 812 -116
rect 814 -156 815 -116
rect 844 -156 845 -116
rect 847 -156 848 -116
rect 269 -379 270 -339
rect 272 -379 273 -339
rect 302 -379 303 -339
rect 305 -379 306 -339
rect 339 -378 340 -338
rect 342 -378 343 -338
rect 378 -374 379 -334
rect 381 -374 382 -334
rect 411 -368 412 -328
rect 414 -368 415 -328
rect 579 -347 580 -307
rect 582 -347 583 -307
rect 612 -341 613 -301
rect 615 -341 616 -301
<< ndcontact >>
rect 252 670 272 674
rect 252 662 272 666
rect 252 584 272 588
rect 797 624 837 628
rect 851 622 855 642
rect 859 622 863 642
rect 797 616 837 620
rect 252 576 272 580
rect 199 556 203 576
rect 207 556 211 576
rect 308 567 312 587
rect 316 567 320 587
rect 341 567 345 587
rect 349 567 353 587
rect 424 574 464 578
rect 478 572 482 592
rect 486 572 490 592
rect 594 595 634 599
rect 648 593 652 613
rect 656 593 660 613
rect 797 605 837 609
rect 797 597 837 601
rect 594 587 634 591
rect 797 586 837 590
rect 424 566 464 570
rect 594 576 634 580
rect 797 578 837 582
rect 594 568 634 572
rect 797 567 837 571
rect 424 555 464 559
rect 594 557 634 561
rect 797 559 837 563
rect 424 547 464 551
rect 594 549 634 553
rect 797 548 837 552
rect 264 532 284 536
rect 424 536 464 540
rect 594 538 634 542
rect 797 540 837 544
rect 424 528 464 532
rect 594 530 634 534
rect 264 524 284 528
rect 264 446 284 450
rect 264 438 284 442
rect 211 418 215 438
rect 219 418 223 438
rect 320 429 324 449
rect 328 429 332 449
rect 353 429 357 449
rect 361 429 365 449
rect 440 432 480 436
rect 494 430 498 450
rect 502 430 506 450
rect 440 424 480 428
rect 610 434 650 438
rect 664 432 668 452
rect 672 432 676 452
rect 610 426 650 430
rect 440 413 480 417
rect 610 415 650 419
rect 440 405 480 409
rect 610 407 650 411
rect 317 394 337 398
rect 317 386 337 390
rect 440 394 480 398
rect 610 396 650 400
rect 440 386 480 390
rect 610 388 650 392
rect 610 378 650 382
rect 686 378 690 398
rect 694 378 698 398
rect 707 378 711 398
rect 715 378 719 398
rect 736 378 740 398
rect 744 378 748 398
rect 769 378 773 398
rect 777 378 781 398
rect 796 378 800 398
rect 804 378 808 398
rect 610 370 650 374
rect 317 308 337 312
rect 818 350 822 370
rect 826 350 830 370
rect 838 350 842 370
rect 846 350 850 370
rect 859 350 863 370
rect 867 350 871 370
rect 888 350 892 370
rect 896 350 900 370
rect 921 350 925 370
rect 929 350 933 370
rect 948 350 952 370
rect 956 350 960 370
rect 317 300 337 304
rect 264 280 268 300
rect 272 280 276 300
rect 373 291 377 311
rect 381 291 385 311
rect 406 291 410 311
rect 414 291 418 311
rect 496 271 536 275
rect 550 269 554 289
rect 558 269 562 289
rect 496 263 536 267
rect 317 256 337 260
rect 317 248 337 252
rect 496 252 536 256
rect 496 244 536 248
rect 593 239 597 259
rect 601 239 605 259
rect 622 239 626 259
rect 630 239 634 259
rect 655 239 659 259
rect 663 239 667 259
rect 682 239 686 259
rect 690 239 694 259
rect 784 261 804 265
rect 496 233 536 237
rect 731 234 735 254
rect 739 234 743 254
rect 784 253 804 257
rect 816 233 820 253
rect 824 233 828 253
rect 840 245 844 265
rect 848 245 852 265
rect 873 245 877 265
rect 881 245 885 265
rect 496 225 536 229
rect 317 170 337 174
rect 317 162 337 166
rect 264 142 268 162
rect 272 142 276 162
rect 373 153 377 173
rect 381 153 385 173
rect 406 153 410 173
rect 414 153 418 173
rect 628 139 648 143
rect 628 131 648 135
rect 264 85 268 105
rect 272 85 276 105
rect 297 85 301 105
rect 305 85 309 105
rect 321 97 325 117
rect 329 97 333 117
rect 345 93 365 97
rect 406 96 410 116
rect 414 96 418 116
rect 450 101 454 121
rect 458 101 462 121
rect 483 101 487 121
rect 491 101 495 121
rect 510 101 514 121
rect 518 101 522 121
rect 345 85 365 89
rect 747 98 767 102
rect 694 71 698 91
rect 702 71 706 91
rect 747 90 767 94
rect 779 70 783 90
rect 787 70 791 90
rect 803 82 807 102
rect 811 82 815 102
rect 836 82 840 102
rect 844 82 848 102
rect 628 53 648 57
rect 628 45 648 49
rect 575 25 579 45
rect 583 25 587 45
rect 625 1 645 5
rect 625 -7 645 -3
rect 264 -49 268 -29
rect 272 -49 276 -29
rect 297 -49 301 -29
rect 305 -49 309 -29
rect 321 -37 325 -17
rect 329 -37 333 -17
rect 345 -41 365 -37
rect 406 -38 410 -18
rect 414 -38 418 -18
rect 345 -49 365 -45
rect 746 -48 766 -44
rect 693 -75 697 -55
rect 701 -75 705 -55
rect 746 -56 766 -52
rect 778 -76 782 -56
rect 786 -76 790 -56
rect 802 -64 806 -44
rect 810 -64 814 -44
rect 835 -64 839 -44
rect 843 -64 847 -44
rect 625 -85 645 -81
rect 625 -93 645 -89
rect 572 -113 576 -93
rect 580 -113 584 -93
rect 628 -137 648 -133
rect 628 -145 648 -141
rect 265 -183 269 -163
rect 273 -183 277 -163
rect 298 -183 302 -163
rect 306 -183 310 -163
rect 322 -171 326 -151
rect 330 -171 334 -151
rect 346 -175 366 -171
rect 407 -172 411 -152
rect 415 -172 419 -152
rect 346 -183 366 -179
rect 751 -182 771 -178
rect 698 -209 702 -189
rect 706 -209 710 -189
rect 751 -190 771 -186
rect 783 -210 787 -190
rect 791 -210 795 -190
rect 807 -198 811 -178
rect 815 -198 819 -178
rect 840 -198 844 -178
rect 848 -198 852 -178
rect 628 -223 648 -219
rect 628 -231 648 -227
rect 575 -251 579 -231
rect 583 -251 587 -231
rect 628 -275 648 -271
rect 628 -283 648 -279
rect 265 -317 269 -297
rect 273 -317 277 -297
rect 298 -317 302 -297
rect 306 -317 310 -297
rect 322 -305 326 -285
rect 330 -305 334 -285
rect 346 -309 366 -305
rect 407 -306 411 -286
rect 415 -306 419 -286
rect 346 -317 366 -313
rect 628 -361 648 -357
rect 628 -369 648 -365
rect 575 -389 579 -369
rect 583 -389 587 -369
<< pdcontact >>
rect 199 598 203 638
rect 207 598 211 638
rect 232 604 236 644
rect 240 604 244 644
rect 308 609 312 649
rect 316 609 320 649
rect 341 609 345 649
rect 349 609 353 649
rect 374 614 378 654
rect 382 614 386 654
rect 407 614 411 654
rect 415 614 419 654
rect 440 614 444 654
rect 448 614 452 654
rect 478 614 482 654
rect 486 614 490 654
rect 511 635 515 675
rect 519 635 523 675
rect 544 635 548 675
rect 552 635 556 675
rect 577 635 581 675
rect 585 635 589 675
rect 610 635 614 675
rect 618 635 622 675
rect 648 635 652 675
rect 656 635 660 675
rect 681 664 685 704
rect 689 664 693 704
rect 714 664 718 704
rect 722 664 726 704
rect 747 664 751 704
rect 755 664 759 704
rect 780 664 784 704
rect 788 664 792 704
rect 813 664 817 704
rect 821 664 825 704
rect 851 664 855 704
rect 859 664 863 704
rect 885 532 925 536
rect 732 527 772 531
rect 885 524 925 528
rect 732 519 772 523
rect 211 460 215 500
rect 219 460 223 500
rect 244 466 248 506
rect 252 466 256 506
rect 320 471 324 511
rect 328 471 332 511
rect 353 471 357 511
rect 361 471 365 511
rect 390 472 394 512
rect 398 472 402 512
rect 423 472 427 512
rect 431 472 435 512
rect 456 472 460 512
rect 464 472 468 512
rect 494 472 498 512
rect 502 472 506 512
rect 527 474 531 514
rect 535 474 539 514
rect 560 474 564 514
rect 568 474 572 514
rect 593 474 597 514
rect 601 474 605 514
rect 626 474 630 514
rect 634 474 638 514
rect 664 474 668 514
rect 672 474 676 514
rect 884 499 924 503
rect 731 493 771 497
rect 884 491 924 495
rect 731 485 771 489
rect 883 465 923 469
rect 731 458 771 462
rect 731 450 771 454
rect 731 425 771 429
rect 731 417 771 421
rect 796 420 800 460
rect 804 420 808 460
rect 883 457 923 461
rect 883 430 923 434
rect 883 422 923 426
rect 883 397 923 401
rect 883 389 923 393
rect 948 392 952 432
rect 956 392 960 432
rect 264 322 268 362
rect 272 322 276 362
rect 297 328 301 368
rect 305 328 309 368
rect 373 333 377 373
rect 381 333 385 373
rect 406 333 410 373
rect 414 333 418 373
rect 617 354 657 358
rect 446 311 450 351
rect 454 311 458 351
rect 479 311 483 351
rect 487 311 491 351
rect 512 311 516 351
rect 520 311 524 351
rect 550 311 554 351
rect 558 311 562 351
rect 617 346 657 350
rect 617 319 657 323
rect 617 311 657 315
rect 617 286 657 290
rect 617 278 657 282
rect 682 281 686 321
rect 690 281 694 321
rect 731 276 735 316
rect 739 276 743 316
rect 764 282 768 322
rect 772 282 776 322
rect 803 286 807 326
rect 811 286 815 326
rect 840 287 844 327
rect 848 287 852 327
rect 873 287 877 327
rect 881 287 885 327
rect 264 184 268 224
rect 272 184 276 224
rect 297 190 301 230
rect 305 190 309 230
rect 373 195 377 235
rect 381 195 385 235
rect 406 195 410 235
rect 414 195 418 235
rect 445 181 485 185
rect 445 173 485 177
rect 445 148 485 152
rect 445 140 485 144
rect 510 143 514 183
rect 518 143 522 183
rect 694 113 698 153
rect 702 113 706 153
rect 727 119 731 159
rect 735 119 739 159
rect 766 123 770 163
rect 774 123 778 163
rect 803 124 807 164
rect 811 124 815 164
rect 836 124 840 164
rect 844 124 848 164
rect 264 23 268 63
rect 272 23 276 63
rect 297 23 301 63
rect 305 23 309 63
rect 334 24 338 64
rect 342 24 346 64
rect 373 28 377 68
rect 381 28 385 68
rect 406 34 410 74
rect 414 34 418 74
rect 575 67 579 107
rect 583 67 587 107
rect 608 73 612 113
rect 616 73 620 113
rect 264 -111 268 -71
rect 272 -111 276 -71
rect 297 -111 301 -71
rect 305 -111 309 -71
rect 334 -110 338 -70
rect 342 -110 346 -70
rect 373 -106 377 -66
rect 381 -106 385 -66
rect 406 -100 410 -60
rect 414 -100 418 -60
rect 572 -71 576 -31
rect 580 -71 584 -31
rect 605 -65 609 -25
rect 613 -65 617 -25
rect 693 -33 697 7
rect 701 -33 705 7
rect 726 -27 730 13
rect 734 -27 738 13
rect 765 -23 769 17
rect 773 -23 777 17
rect 802 -22 806 18
rect 810 -22 814 18
rect 835 -22 839 18
rect 843 -22 847 18
rect 265 -245 269 -205
rect 273 -245 277 -205
rect 298 -245 302 -205
rect 306 -245 310 -205
rect 335 -244 339 -204
rect 343 -244 347 -204
rect 374 -240 378 -200
rect 382 -240 386 -200
rect 407 -234 411 -194
rect 415 -234 419 -194
rect 575 -209 579 -169
rect 583 -209 587 -169
rect 608 -203 612 -163
rect 616 -203 620 -163
rect 698 -167 702 -127
rect 706 -167 710 -127
rect 731 -161 735 -121
rect 739 -161 743 -121
rect 770 -157 774 -117
rect 778 -157 782 -117
rect 807 -156 811 -116
rect 815 -156 819 -116
rect 840 -156 844 -116
rect 848 -156 852 -116
rect 265 -379 269 -339
rect 273 -379 277 -339
rect 298 -379 302 -339
rect 306 -379 310 -339
rect 335 -378 339 -338
rect 343 -378 347 -338
rect 374 -374 378 -334
rect 382 -374 386 -334
rect 407 -368 411 -328
rect 415 -368 419 -328
rect 575 -347 579 -307
rect 583 -347 587 -307
rect 608 -341 612 -301
rect 616 -341 620 -301
<< polysilicon >>
rect 686 704 688 707
rect 719 704 721 707
rect 752 704 754 707
rect 785 704 787 707
rect 818 704 820 707
rect 856 704 858 707
rect 516 675 518 678
rect 549 675 551 678
rect 582 675 584 678
rect 615 675 617 678
rect 653 675 655 678
rect 249 667 252 669
rect 272 667 275 669
rect 379 654 381 657
rect 412 654 414 657
rect 445 654 447 657
rect 483 654 485 657
rect 313 649 315 652
rect 346 649 348 652
rect 237 644 239 647
rect 204 638 206 641
rect 686 651 688 664
rect 719 651 721 664
rect 752 651 754 664
rect 785 651 787 664
rect 818 651 820 664
rect 856 642 858 664
rect 516 622 518 635
rect 549 622 551 635
rect 582 622 584 635
rect 615 622 617 635
rect 204 576 206 598
rect 237 592 239 604
rect 313 587 315 609
rect 346 587 348 609
rect 379 601 381 614
rect 412 601 414 614
rect 445 601 447 614
rect 483 592 485 614
rect 653 613 655 635
rect 794 621 797 623
rect 837 621 840 623
rect 856 619 858 622
rect 244 581 252 583
rect 272 581 275 583
rect 421 571 424 573
rect 464 571 467 573
rect 591 592 594 594
rect 634 592 637 594
rect 794 602 797 604
rect 837 602 840 604
rect 653 590 655 593
rect 794 583 797 585
rect 837 583 840 585
rect 313 564 315 567
rect 346 564 348 567
rect 483 569 485 572
rect 591 573 594 575
rect 634 573 637 575
rect 794 564 797 566
rect 837 564 840 566
rect 204 553 206 556
rect 421 552 424 554
rect 464 552 467 554
rect 591 554 594 556
rect 634 554 637 556
rect 794 545 797 547
rect 837 545 840 547
rect 421 533 424 535
rect 464 533 467 535
rect 591 535 594 537
rect 634 535 637 537
rect 261 529 264 531
rect 284 529 287 531
rect 882 529 885 531
rect 925 529 936 531
rect 729 524 732 526
rect 772 524 783 526
rect 325 511 327 514
rect 358 511 360 514
rect 395 512 397 515
rect 428 512 430 515
rect 461 512 463 515
rect 499 512 501 515
rect 532 514 534 517
rect 565 514 567 517
rect 598 514 600 517
rect 631 514 633 517
rect 669 514 671 517
rect 249 506 251 509
rect 216 500 218 503
rect 881 496 884 498
rect 924 496 935 498
rect 728 490 731 492
rect 771 490 782 492
rect 216 438 218 460
rect 249 454 251 466
rect 325 449 327 471
rect 358 449 360 471
rect 395 459 397 472
rect 428 459 430 472
rect 461 459 463 472
rect 499 450 501 472
rect 532 461 534 474
rect 565 461 567 474
rect 598 461 600 474
rect 631 461 633 474
rect 669 452 671 474
rect 801 460 803 463
rect 880 462 883 464
rect 923 462 934 464
rect 728 455 731 457
rect 771 455 782 457
rect 256 443 264 445
rect 284 443 287 445
rect 325 426 327 429
rect 358 426 360 429
rect 437 429 440 431
rect 480 429 483 431
rect 499 427 501 430
rect 607 431 610 433
rect 650 431 653 433
rect 669 429 671 432
rect 728 422 731 424
rect 771 422 777 424
rect 216 415 218 418
rect 437 410 440 412
rect 480 410 483 412
rect 775 418 777 422
rect 953 432 955 435
rect 880 427 883 429
rect 923 427 934 429
rect 607 412 610 414
rect 650 412 653 414
rect 314 391 317 393
rect 337 391 340 393
rect 437 391 440 393
rect 480 391 483 393
rect 691 398 693 401
rect 712 398 714 401
rect 741 398 743 401
rect 774 398 776 401
rect 801 398 803 420
rect 607 393 610 395
rect 650 393 653 395
rect 378 373 380 376
rect 411 373 413 376
rect 880 394 883 396
rect 923 394 929 396
rect 927 390 929 394
rect 607 375 610 377
rect 650 375 653 377
rect 691 375 693 378
rect 712 375 714 378
rect 741 375 743 378
rect 774 375 776 378
rect 801 375 803 378
rect 302 368 304 371
rect 269 362 271 365
rect 823 370 825 373
rect 843 370 845 373
rect 864 370 866 373
rect 893 370 895 373
rect 926 370 928 373
rect 953 370 955 392
rect 451 351 453 354
rect 484 351 486 354
rect 517 351 519 354
rect 555 351 557 354
rect 269 300 271 322
rect 302 316 304 328
rect 378 311 380 333
rect 411 311 413 333
rect 614 351 617 353
rect 657 351 668 353
rect 823 347 825 350
rect 843 347 845 350
rect 864 347 866 350
rect 893 347 895 350
rect 926 347 928 350
rect 953 347 955 350
rect 808 326 810 329
rect 845 327 847 330
rect 878 327 880 330
rect 687 321 689 324
rect 769 322 771 325
rect 614 316 617 318
rect 657 316 668 318
rect 309 305 317 307
rect 337 305 340 307
rect 451 298 453 311
rect 484 298 486 311
rect 517 298 519 311
rect 378 288 380 291
rect 411 288 413 291
rect 555 289 557 311
rect 269 277 271 280
rect 493 268 496 270
rect 536 268 539 270
rect 614 283 617 285
rect 657 283 663 285
rect 661 279 663 283
rect 736 316 738 319
rect 555 266 557 269
rect 598 259 600 262
rect 627 259 629 262
rect 660 259 662 262
rect 687 259 689 281
rect 808 283 810 286
rect 769 276 771 282
rect 314 253 317 255
rect 337 253 340 255
rect 493 249 496 251
rect 536 249 539 251
rect 736 254 738 276
rect 845 265 847 287
rect 878 265 880 287
rect 776 258 784 260
rect 804 258 807 260
rect 378 235 380 238
rect 411 235 413 238
rect 302 230 304 233
rect 269 224 271 227
rect 598 236 600 239
rect 627 236 629 239
rect 660 236 662 239
rect 687 236 689 239
rect 821 253 823 257
rect 493 230 496 232
rect 536 230 539 232
rect 736 231 738 234
rect 845 242 847 245
rect 878 242 880 245
rect 821 230 823 233
rect 269 162 271 184
rect 302 178 304 190
rect 378 173 380 195
rect 411 173 413 195
rect 515 183 517 186
rect 442 178 445 180
rect 485 178 496 180
rect 309 167 317 169
rect 337 167 340 169
rect 378 150 380 153
rect 411 150 413 153
rect 442 145 445 147
rect 485 145 491 147
rect 269 139 271 142
rect 489 141 491 145
rect 771 163 773 166
rect 808 164 810 167
rect 841 164 843 167
rect 732 159 734 162
rect 699 153 701 156
rect 455 121 457 124
rect 488 121 490 124
rect 515 121 517 143
rect 625 136 628 138
rect 648 136 651 138
rect 326 117 328 120
rect 269 105 271 108
rect 302 105 304 108
rect 411 116 413 119
rect 326 93 328 97
rect 613 113 615 116
rect 771 120 773 123
rect 732 113 734 119
rect 580 107 582 110
rect 455 98 457 101
rect 488 98 490 101
rect 515 98 517 101
rect 342 90 345 92
rect 365 90 373 92
rect 269 63 271 85
rect 302 63 304 85
rect 411 74 413 96
rect 378 68 380 74
rect 339 64 341 67
rect 699 91 701 113
rect 808 102 810 124
rect 841 102 843 124
rect 739 95 747 97
rect 767 95 770 97
rect 580 45 582 67
rect 613 61 615 73
rect 784 90 786 94
rect 699 68 701 71
rect 808 79 810 82
rect 841 79 843 82
rect 784 67 786 70
rect 620 50 628 52
rect 648 50 651 52
rect 411 31 413 34
rect 378 25 380 28
rect 269 20 271 23
rect 302 20 304 23
rect 339 21 341 24
rect 580 22 582 25
rect 770 17 772 20
rect 807 18 809 21
rect 840 18 842 21
rect 731 13 733 16
rect 698 7 700 10
rect 622 -2 625 0
rect 645 -2 648 0
rect 326 -17 328 -14
rect 269 -29 271 -26
rect 302 -29 304 -26
rect 411 -18 413 -15
rect 326 -41 328 -37
rect 610 -25 612 -22
rect 577 -31 579 -28
rect 342 -44 345 -42
rect 365 -44 373 -42
rect 269 -71 271 -49
rect 302 -71 304 -49
rect 411 -60 413 -38
rect 378 -66 380 -60
rect 339 -70 341 -67
rect 770 -26 772 -23
rect 731 -33 733 -27
rect 698 -55 700 -33
rect 807 -44 809 -22
rect 840 -44 842 -22
rect 738 -51 746 -49
rect 766 -51 769 -49
rect 577 -93 579 -71
rect 610 -77 612 -65
rect 783 -56 785 -52
rect 698 -78 700 -75
rect 807 -67 809 -64
rect 840 -67 842 -64
rect 783 -79 785 -76
rect 617 -88 625 -86
rect 645 -88 648 -86
rect 411 -103 413 -100
rect 378 -109 380 -106
rect 269 -114 271 -111
rect 302 -114 304 -111
rect 339 -113 341 -110
rect 577 -116 579 -113
rect 775 -117 777 -114
rect 812 -116 814 -113
rect 845 -116 847 -113
rect 736 -121 738 -118
rect 703 -127 705 -124
rect 625 -140 628 -138
rect 648 -140 651 -138
rect 327 -151 329 -148
rect 270 -163 272 -160
rect 303 -163 305 -160
rect 412 -152 414 -149
rect 327 -175 329 -171
rect 613 -163 615 -160
rect 580 -169 582 -166
rect 343 -178 346 -176
rect 366 -178 374 -176
rect 270 -205 272 -183
rect 303 -205 305 -183
rect 412 -194 414 -172
rect 379 -200 381 -194
rect 340 -204 342 -201
rect 775 -160 777 -157
rect 736 -167 738 -161
rect 703 -189 705 -167
rect 812 -178 814 -156
rect 845 -178 847 -156
rect 743 -185 751 -183
rect 771 -185 774 -183
rect 580 -231 582 -209
rect 613 -215 615 -203
rect 788 -190 790 -186
rect 703 -212 705 -209
rect 812 -201 814 -198
rect 845 -201 847 -198
rect 788 -213 790 -210
rect 620 -226 628 -224
rect 648 -226 651 -224
rect 412 -237 414 -234
rect 379 -243 381 -240
rect 270 -248 272 -245
rect 303 -248 305 -245
rect 340 -247 342 -244
rect 580 -254 582 -251
rect 625 -278 628 -276
rect 648 -278 651 -276
rect 327 -285 329 -282
rect 270 -297 272 -294
rect 303 -297 305 -294
rect 412 -286 414 -283
rect 327 -309 329 -305
rect 613 -301 615 -298
rect 343 -312 346 -310
rect 366 -312 374 -310
rect 270 -339 272 -317
rect 303 -339 305 -317
rect 412 -328 414 -306
rect 580 -307 582 -304
rect 379 -334 381 -328
rect 340 -338 342 -335
rect 412 -371 414 -368
rect 580 -369 582 -347
rect 613 -353 615 -341
rect 620 -364 628 -362
rect 648 -364 651 -362
rect 379 -377 381 -374
rect 270 -382 272 -379
rect 303 -382 305 -379
rect 340 -381 342 -378
rect 580 -392 582 -389
<< polycontact >>
rect 245 666 249 670
rect 685 647 689 651
rect 718 647 722 651
rect 751 647 755 651
rect 784 647 788 651
rect 817 647 821 651
rect 852 646 856 650
rect 515 618 519 622
rect 548 618 552 622
rect 581 618 585 622
rect 614 618 618 622
rect 649 617 653 621
rect 200 580 204 584
rect 236 588 240 592
rect 309 591 313 595
rect 342 591 346 595
rect 378 597 382 601
rect 411 597 415 601
rect 444 597 448 601
rect 479 596 483 600
rect 788 619 794 625
rect 240 580 244 584
rect 415 569 421 575
rect 585 590 591 596
rect 788 600 794 606
rect 788 581 794 587
rect 585 571 591 577
rect 788 562 794 568
rect 415 550 421 556
rect 585 552 591 558
rect 788 543 794 549
rect 257 528 261 532
rect 415 531 421 537
rect 585 533 591 539
rect 878 528 882 532
rect 725 523 729 527
rect 877 495 881 499
rect 724 489 728 493
rect 212 442 216 446
rect 248 450 252 454
rect 321 453 325 457
rect 354 453 358 457
rect 394 455 398 459
rect 427 455 431 459
rect 460 455 464 459
rect 495 454 499 458
rect 531 457 535 461
rect 564 457 568 461
rect 597 457 601 461
rect 630 457 634 461
rect 665 456 669 460
rect 876 461 880 465
rect 724 454 728 458
rect 252 442 256 446
rect 431 427 437 433
rect 601 429 607 435
rect 431 408 437 414
rect 601 410 607 416
rect 876 426 880 430
rect 774 414 778 418
rect 690 401 694 405
rect 711 401 715 405
rect 740 401 744 405
rect 774 401 778 405
rect 797 402 801 406
rect 310 390 314 394
rect 431 389 437 395
rect 601 391 607 397
rect 601 373 607 379
rect 926 386 930 390
rect 822 373 826 377
rect 842 373 846 377
rect 863 373 867 377
rect 892 373 896 377
rect 926 373 930 377
rect 949 374 953 378
rect 265 304 269 308
rect 301 312 305 316
rect 374 315 378 319
rect 407 315 411 319
rect 610 350 614 354
rect 768 325 772 329
rect 610 315 614 319
rect 305 304 309 308
rect 450 294 454 298
rect 483 294 487 298
rect 516 294 520 298
rect 551 293 555 297
rect 487 266 493 272
rect 660 275 664 279
rect 597 262 601 266
rect 626 262 630 266
rect 660 262 664 266
rect 683 263 687 267
rect 806 278 812 283
rect 310 252 314 256
rect 487 247 493 253
rect 732 258 736 262
rect 841 269 845 273
rect 874 269 878 273
rect 772 257 776 261
rect 819 257 825 262
rect 487 228 493 234
rect 265 166 269 170
rect 301 174 305 178
rect 374 177 378 181
rect 407 177 411 181
rect 438 177 442 181
rect 305 166 309 170
rect 731 162 735 166
rect 488 137 492 141
rect 454 124 458 128
rect 488 124 492 128
rect 511 125 515 129
rect 621 135 625 139
rect 769 115 775 120
rect 324 88 330 93
rect 373 89 377 93
rect 271 77 275 81
rect 304 77 308 81
rect 413 88 417 92
rect 337 67 343 72
rect 695 95 699 99
rect 804 106 808 110
rect 837 106 841 110
rect 735 94 739 98
rect 782 94 788 99
rect 576 49 580 53
rect 612 57 616 61
rect 616 49 620 53
rect 377 21 381 25
rect 730 16 734 20
rect 618 -3 622 1
rect 324 -46 330 -41
rect 373 -45 377 -41
rect 271 -57 275 -53
rect 304 -57 308 -53
rect 413 -46 417 -42
rect 337 -67 343 -62
rect 768 -31 774 -26
rect 694 -51 698 -47
rect 803 -40 807 -36
rect 836 -40 840 -36
rect 734 -52 738 -48
rect 781 -52 787 -47
rect 573 -89 577 -85
rect 609 -81 613 -77
rect 613 -89 617 -85
rect 377 -113 381 -109
rect 735 -118 739 -114
rect 621 -141 625 -137
rect 325 -180 331 -175
rect 374 -179 378 -175
rect 272 -191 276 -187
rect 305 -191 309 -187
rect 414 -180 418 -176
rect 338 -201 344 -196
rect 773 -165 779 -160
rect 699 -185 703 -181
rect 808 -174 812 -170
rect 841 -174 845 -170
rect 739 -186 743 -182
rect 786 -186 792 -181
rect 576 -227 580 -223
rect 612 -219 616 -215
rect 616 -227 620 -223
rect 378 -247 382 -243
rect 621 -279 625 -275
rect 325 -314 331 -309
rect 374 -313 378 -309
rect 272 -325 276 -321
rect 305 -325 309 -321
rect 414 -314 418 -310
rect 338 -335 344 -330
rect 576 -365 580 -361
rect 612 -357 616 -353
rect 616 -365 620 -361
rect 378 -381 382 -377
<< metal1 >>
rect 675 714 869 717
rect 675 710 699 714
rect 708 710 732 714
rect 741 710 765 714
rect 774 710 798 714
rect 807 710 831 714
rect 845 710 869 714
rect 681 704 685 710
rect 714 704 718 710
rect 747 704 751 710
rect 780 704 784 710
rect 813 704 817 710
rect 851 704 855 710
rect 505 685 666 688
rect 505 681 529 685
rect 538 681 562 685
rect 571 681 595 685
rect 604 681 628 685
rect 642 681 666 685
rect 511 675 515 681
rect 544 675 548 681
rect 577 675 581 681
rect 610 675 614 681
rect 648 675 652 681
rect 272 670 285 674
rect 185 666 245 670
rect 185 584 190 666
rect 268 653 272 662
rect 193 644 217 651
rect 226 650 272 653
rect 232 644 236 650
rect 199 638 203 644
rect 207 584 211 598
rect 240 599 244 604
rect 279 599 285 670
rect 368 664 496 667
rect 302 655 359 662
rect 368 660 392 664
rect 401 660 425 664
rect 434 660 458 664
rect 472 660 496 664
rect 308 649 312 655
rect 341 649 345 655
rect 374 654 378 660
rect 407 654 411 660
rect 440 654 444 660
rect 478 654 482 660
rect 689 654 693 664
rect 722 654 726 664
rect 755 654 759 664
rect 788 654 792 664
rect 821 654 825 664
rect 519 625 523 635
rect 552 625 556 635
rect 585 625 589 635
rect 618 625 622 635
rect 240 596 285 599
rect 240 595 302 596
rect 316 595 320 609
rect 349 595 353 609
rect 382 604 386 614
rect 415 604 419 614
rect 448 604 452 614
rect 236 584 240 588
rect 272 584 276 595
rect 282 591 309 595
rect 316 591 342 595
rect 349 591 361 595
rect 316 587 320 591
rect 349 587 353 591
rect 185 580 200 584
rect 207 580 240 584
rect 207 576 211 580
rect 199 547 203 556
rect 268 547 272 576
rect 308 547 312 567
rect 341 547 345 567
rect 193 539 360 547
rect 378 537 382 597
rect 401 597 411 601
rect 486 600 490 614
rect 401 556 405 597
rect 444 592 448 597
rect 415 589 448 592
rect 460 596 479 600
rect 486 596 501 600
rect 415 575 421 589
rect 460 578 464 596
rect 486 592 490 596
rect 478 570 482 572
rect 460 559 464 566
rect 401 550 415 556
rect 472 567 482 570
rect 460 540 464 547
rect 284 532 297 536
rect 197 528 257 532
rect 197 446 202 528
rect 280 515 284 524
rect 205 506 229 513
rect 238 512 284 515
rect 244 506 248 512
rect 211 500 215 506
rect 219 446 223 460
rect 252 461 256 466
rect 291 461 297 532
rect 378 531 415 537
rect 472 532 476 567
rect 515 539 519 618
rect 548 558 552 618
rect 571 618 581 622
rect 656 621 660 635
rect 571 577 575 618
rect 614 613 618 618
rect 585 610 618 613
rect 630 617 649 621
rect 656 617 671 621
rect 585 596 591 610
rect 630 599 634 617
rect 656 613 660 617
rect 648 591 652 593
rect 630 580 634 587
rect 571 571 585 577
rect 642 588 652 591
rect 630 561 634 568
rect 548 552 585 558
rect 630 542 634 549
rect 515 533 585 539
rect 642 534 646 588
rect 685 549 689 647
rect 718 568 722 647
rect 751 587 755 647
rect 774 647 784 651
rect 859 650 863 664
rect 774 606 778 647
rect 817 642 821 647
rect 788 639 821 642
rect 833 646 852 650
rect 859 646 874 650
rect 788 625 794 639
rect 833 628 837 646
rect 859 642 863 646
rect 851 620 855 622
rect 833 609 837 616
rect 774 600 788 606
rect 845 617 855 620
rect 833 590 837 597
rect 751 581 788 587
rect 833 571 837 578
rect 718 562 788 568
rect 833 552 837 559
rect 685 543 788 549
rect 845 544 849 617
rect 837 540 849 544
rect 464 528 476 532
rect 634 530 646 534
rect 925 532 947 536
rect 772 527 795 531
rect 314 517 371 524
rect 384 522 512 525
rect 384 518 408 522
rect 417 518 441 522
rect 450 518 474 522
rect 488 518 512 522
rect 521 524 682 527
rect 521 520 545 524
rect 554 520 578 524
rect 587 520 611 524
rect 620 520 644 524
rect 658 520 682 524
rect 690 523 725 527
rect 320 511 324 517
rect 353 511 357 517
rect 390 512 394 518
rect 423 512 427 518
rect 456 512 460 518
rect 494 512 498 518
rect 527 514 531 520
rect 560 514 564 520
rect 593 514 597 520
rect 626 514 630 520
rect 664 514 668 520
rect 252 458 297 461
rect 252 457 314 458
rect 328 457 332 471
rect 361 457 365 471
rect 398 462 402 472
rect 431 462 435 472
rect 464 462 468 472
rect 248 446 252 450
rect 284 446 288 457
rect 294 453 321 457
rect 328 453 354 457
rect 361 453 373 457
rect 328 449 332 453
rect 361 449 365 453
rect 197 442 212 446
rect 219 442 252 446
rect 219 438 223 442
rect 211 409 215 418
rect 280 409 284 438
rect 320 409 324 429
rect 353 409 357 429
rect 205 401 372 409
rect 337 394 350 398
rect 250 390 310 394
rect 250 308 255 390
rect 333 377 337 386
rect 258 368 282 375
rect 291 374 337 377
rect 297 368 301 374
rect 264 362 268 368
rect 272 308 276 322
rect 305 323 309 328
rect 344 323 350 394
rect 394 395 398 455
rect 417 455 427 459
rect 502 458 506 472
rect 535 464 539 474
rect 568 464 572 474
rect 601 464 605 474
rect 634 464 638 474
rect 417 414 421 455
rect 460 450 464 455
rect 431 447 464 450
rect 476 454 495 458
rect 502 454 517 458
rect 431 433 437 447
rect 476 436 480 454
rect 502 450 506 454
rect 494 428 498 430
rect 476 417 480 424
rect 417 408 431 414
rect 488 425 498 428
rect 476 398 480 405
rect 394 389 431 395
rect 488 390 492 425
rect 480 386 492 390
rect 367 379 424 386
rect 531 379 535 457
rect 564 397 568 457
rect 587 457 597 461
rect 672 460 676 474
rect 587 416 591 457
rect 630 452 634 457
rect 601 449 634 452
rect 646 456 665 460
rect 672 456 687 460
rect 601 435 607 449
rect 646 438 650 456
rect 672 452 676 456
rect 664 430 668 432
rect 646 419 650 426
rect 587 410 601 416
rect 658 427 668 430
rect 646 400 650 407
rect 564 391 601 397
rect 646 382 650 388
rect 373 373 377 379
rect 406 373 410 379
rect 531 373 601 379
rect 658 374 662 427
rect 690 405 694 523
rect 767 497 772 519
rect 771 493 772 497
rect 711 489 724 493
rect 711 405 715 489
rect 766 462 771 485
rect 790 473 795 527
rect 822 528 878 532
rect 790 466 814 473
rect 796 460 800 466
rect 731 444 735 450
rect 723 440 735 444
rect 723 421 727 440
rect 771 425 787 429
rect 723 417 731 421
rect 774 405 778 414
rect 782 406 787 425
rect 804 406 808 420
rect 782 402 797 406
rect 804 402 819 406
rect 650 370 662 374
rect 787 394 791 402
rect 804 398 808 402
rect 686 374 690 378
rect 707 374 711 378
rect 736 374 740 378
rect 769 374 773 378
rect 796 374 800 378
rect 686 371 800 374
rect 822 377 826 528
rect 920 503 925 524
rect 924 499 925 503
rect 842 495 877 499
rect 842 377 846 495
rect 919 469 924 491
rect 923 465 924 469
rect 863 461 876 465
rect 863 377 867 461
rect 918 434 923 457
rect 942 445 947 532
rect 942 438 966 445
rect 948 432 952 438
rect 883 416 887 422
rect 875 412 887 416
rect 875 393 879 412
rect 923 397 939 401
rect 875 389 883 393
rect 926 377 930 386
rect 934 378 939 397
rect 956 378 960 392
rect 934 374 949 378
rect 956 374 971 378
rect 440 361 568 364
rect 440 357 464 361
rect 473 357 497 361
rect 506 357 530 361
rect 544 357 568 361
rect 305 320 350 323
rect 305 319 367 320
rect 381 319 385 333
rect 414 319 418 333
rect 446 351 450 357
rect 479 351 483 357
rect 512 351 516 357
rect 550 351 554 357
rect 657 354 681 358
rect 301 308 305 312
rect 337 308 341 319
rect 347 315 374 319
rect 381 315 407 319
rect 414 315 426 319
rect 381 311 385 315
rect 414 311 418 315
rect 209 304 265 308
rect 272 304 305 308
rect 209 -53 216 304
rect 272 300 276 304
rect 264 271 268 280
rect 333 271 337 300
rect 454 301 458 311
rect 487 301 491 311
rect 520 301 524 311
rect 373 271 377 291
rect 406 271 410 291
rect 257 263 424 271
rect 337 256 350 260
rect 250 252 310 256
rect 250 170 255 252
rect 333 239 337 248
rect 258 230 282 237
rect 291 236 337 239
rect 297 230 301 236
rect 264 224 268 230
rect 272 170 276 184
rect 305 185 309 190
rect 344 185 350 256
rect 367 241 424 248
rect 373 235 377 241
rect 406 235 410 241
rect 450 234 454 294
rect 473 294 483 298
rect 558 297 562 311
rect 597 350 610 354
rect 473 253 477 294
rect 516 289 520 294
rect 487 286 520 289
rect 532 293 551 297
rect 558 293 573 297
rect 487 272 493 286
rect 532 275 536 293
rect 558 289 562 293
rect 550 267 554 269
rect 532 256 536 263
rect 473 247 487 253
rect 544 264 554 267
rect 597 266 601 350
rect 652 323 657 346
rect 676 334 681 354
rect 939 366 943 374
rect 956 370 960 374
rect 717 344 807 348
rect 676 327 700 334
rect 682 321 686 327
rect 617 305 621 311
rect 609 301 621 305
rect 609 282 613 301
rect 657 286 673 290
rect 609 278 617 282
rect 660 266 664 275
rect 532 237 536 244
rect 450 228 487 234
rect 544 229 548 264
rect 668 267 673 286
rect 690 267 694 281
rect 668 263 683 267
rect 690 263 705 267
rect 673 255 677 263
rect 690 259 694 263
rect 717 262 722 344
rect 768 329 772 344
rect 725 322 749 329
rect 803 326 807 344
rect 818 346 822 350
rect 838 346 842 350
rect 859 346 863 350
rect 888 346 892 350
rect 921 346 925 350
rect 948 346 952 350
rect 818 343 952 346
rect 834 333 891 340
rect 840 327 844 333
rect 873 327 877 333
rect 731 316 735 322
rect 739 262 743 276
rect 717 258 732 262
rect 739 258 754 262
rect 739 254 743 258
rect 593 235 597 239
rect 622 235 626 239
rect 655 235 659 239
rect 682 235 686 239
rect 593 232 686 235
rect 749 248 754 258
rect 764 261 768 282
rect 815 286 833 290
rect 772 273 776 282
rect 829 273 833 286
rect 848 273 852 287
rect 881 273 885 287
rect 772 269 841 273
rect 848 269 874 273
rect 881 269 893 273
rect 804 261 808 269
rect 764 257 772 261
rect 784 248 788 253
rect 749 244 788 248
rect 536 225 548 229
rect 731 225 735 234
rect 831 250 835 269
rect 848 265 852 269
rect 881 265 885 269
rect 828 247 835 250
rect 816 225 820 233
rect 840 225 844 245
rect 873 225 877 245
rect 725 217 892 225
rect 305 182 350 185
rect 305 181 367 182
rect 381 181 385 195
rect 414 181 418 195
rect 480 191 528 196
rect 480 185 485 191
rect 504 189 528 191
rect 510 183 514 189
rect 301 170 305 174
rect 337 170 341 181
rect 347 177 374 181
rect 381 177 407 181
rect 414 177 438 181
rect 381 173 385 177
rect 414 173 418 177
rect 238 166 265 170
rect 272 166 305 170
rect 238 81 243 166
rect 272 162 276 166
rect 264 133 268 142
rect 333 133 337 162
rect 373 133 377 153
rect 406 133 410 153
rect 257 125 424 133
rect 427 128 431 177
rect 445 167 449 173
rect 437 163 449 167
rect 437 144 441 163
rect 485 148 501 152
rect 437 140 445 144
rect 488 128 492 137
rect 272 105 276 125
rect 305 105 309 125
rect 329 117 333 125
rect 314 100 321 103
rect 264 81 268 85
rect 297 81 301 85
rect 314 81 318 100
rect 414 116 418 125
rect 427 124 454 128
rect 496 129 501 148
rect 680 181 770 185
rect 518 129 522 143
rect 648 139 661 143
rect 561 135 621 139
rect 496 125 511 129
rect 518 125 533 129
rect 361 102 400 106
rect 361 97 365 102
rect 377 89 385 93
rect 341 81 345 89
rect 238 77 268 81
rect 275 77 301 81
rect 308 77 377 81
rect 264 63 268 77
rect 297 63 301 77
rect 316 64 320 77
rect 373 68 377 77
rect 316 60 334 64
rect 381 68 385 89
rect 395 92 400 102
rect 501 117 505 125
rect 518 121 522 125
rect 450 97 454 101
rect 483 97 487 101
rect 510 97 514 101
rect 406 92 410 96
rect 448 94 514 97
rect 395 88 410 92
rect 417 88 432 92
rect 406 74 410 88
rect 414 28 418 34
rect 427 38 432 88
rect 561 53 566 135
rect 644 122 648 131
rect 569 113 593 120
rect 602 119 648 122
rect 608 113 612 119
rect 575 107 579 113
rect 583 53 587 67
rect 616 68 620 73
rect 655 72 661 139
rect 680 99 685 181
rect 731 166 735 181
rect 688 159 712 166
rect 766 163 770 181
rect 797 170 854 177
rect 803 164 807 170
rect 836 164 840 170
rect 694 153 698 159
rect 702 99 706 113
rect 680 95 695 99
rect 702 95 717 99
rect 702 91 706 95
rect 655 68 669 72
rect 616 64 669 68
rect 712 85 717 95
rect 727 98 731 119
rect 778 123 796 127
rect 735 110 739 119
rect 792 110 796 123
rect 811 110 815 124
rect 844 110 848 124
rect 735 106 804 110
rect 811 106 837 110
rect 844 106 856 110
rect 767 98 771 106
rect 727 94 735 98
rect 747 85 751 90
rect 712 81 751 85
rect 612 53 616 57
rect 648 53 652 64
rect 694 62 698 71
rect 794 87 798 106
rect 811 102 815 106
rect 844 102 848 106
rect 791 84 798 87
rect 779 62 783 70
rect 803 62 807 82
rect 836 62 840 82
rect 688 54 855 62
rect 561 49 576 53
rect 583 49 616 53
rect 583 45 587 49
rect 427 30 518 38
rect 272 17 276 23
rect 305 17 309 23
rect 258 10 315 17
rect 342 6 346 24
rect 400 21 424 28
rect 377 6 381 21
rect 427 6 432 30
rect 470 25 518 30
rect 470 9 518 22
rect 575 16 579 25
rect 644 16 648 45
rect 679 35 769 39
rect 569 8 662 16
rect 342 2 432 6
rect 645 1 658 5
rect 257 -9 424 -1
rect 558 -3 618 1
rect 272 -29 276 -9
rect 305 -29 309 -9
rect 329 -17 333 -9
rect 314 -34 321 -31
rect 264 -53 268 -49
rect 297 -53 301 -49
rect 314 -53 318 -34
rect 414 -18 418 -9
rect 361 -32 400 -28
rect 361 -37 365 -32
rect 377 -45 385 -41
rect 341 -53 345 -45
rect 209 -57 268 -53
rect 275 -57 301 -53
rect 308 -57 377 -53
rect 264 -71 268 -57
rect 297 -71 301 -57
rect 316 -70 320 -57
rect 373 -66 377 -57
rect 316 -74 334 -70
rect 381 -66 385 -45
rect 395 -42 400 -32
rect 406 -42 410 -38
rect 395 -46 410 -42
rect 417 -46 432 -42
rect 406 -60 410 -46
rect 414 -106 418 -100
rect 427 -101 432 -46
rect 558 -85 563 -3
rect 641 -16 645 -7
rect 566 -25 590 -18
rect 599 -19 645 -16
rect 605 -25 609 -19
rect 572 -31 576 -25
rect 580 -85 584 -71
rect 613 -70 617 -65
rect 652 -70 658 1
rect 679 -47 684 35
rect 730 20 734 35
rect 687 13 711 20
rect 765 17 769 35
rect 796 24 853 31
rect 802 18 806 24
rect 835 18 839 24
rect 693 7 697 13
rect 701 -47 705 -33
rect 679 -51 694 -47
rect 701 -51 716 -47
rect 701 -55 705 -51
rect 613 -73 658 -70
rect 613 -74 664 -73
rect 609 -85 613 -81
rect 645 -85 649 -74
rect 655 -78 664 -74
rect 711 -61 716 -51
rect 726 -48 730 -27
rect 777 -23 795 -19
rect 734 -36 738 -27
rect 791 -36 795 -23
rect 810 -36 814 -22
rect 843 -36 847 -22
rect 734 -40 803 -36
rect 810 -40 836 -36
rect 843 -40 855 -36
rect 766 -48 770 -40
rect 726 -52 734 -48
rect 746 -61 750 -56
rect 711 -65 750 -61
rect 693 -84 697 -75
rect 793 -59 797 -40
rect 810 -44 814 -40
rect 843 -44 847 -40
rect 790 -62 797 -59
rect 778 -84 782 -76
rect 802 -84 806 -64
rect 835 -84 839 -64
rect 558 -89 573 -85
rect 580 -89 613 -85
rect 580 -93 584 -89
rect 687 -92 854 -84
rect 470 -101 518 -99
rect 272 -117 276 -111
rect 305 -117 309 -111
rect 258 -124 315 -117
rect 342 -128 346 -110
rect 400 -113 424 -106
rect 427 -107 518 -101
rect 377 -128 381 -113
rect 427 -128 432 -107
rect 470 -112 518 -107
rect 470 -127 518 -115
rect 572 -122 576 -113
rect 641 -122 645 -93
rect 684 -99 774 -95
rect 342 -132 432 -128
rect 566 -130 664 -122
rect 258 -143 425 -135
rect 648 -137 661 -133
rect 561 -141 621 -137
rect 273 -163 277 -143
rect 306 -163 310 -143
rect 330 -151 334 -143
rect 315 -168 322 -165
rect 265 -187 269 -183
rect 298 -187 302 -183
rect 315 -187 319 -168
rect 415 -152 419 -143
rect 362 -166 401 -162
rect 362 -171 366 -166
rect 378 -179 386 -175
rect 342 -187 346 -179
rect 257 -191 269 -187
rect 276 -191 302 -187
rect 309 -191 378 -187
rect 265 -205 269 -191
rect 298 -205 302 -191
rect 317 -204 321 -191
rect 374 -200 378 -191
rect 317 -208 335 -204
rect 382 -200 386 -179
rect 396 -176 401 -166
rect 407 -176 411 -172
rect 396 -180 411 -176
rect 418 -180 433 -176
rect 407 -194 411 -180
rect 415 -240 419 -234
rect 428 -240 433 -180
rect 561 -223 566 -141
rect 644 -154 648 -145
rect 569 -163 593 -156
rect 602 -157 648 -154
rect 608 -163 612 -157
rect 575 -169 579 -163
rect 583 -223 587 -209
rect 616 -208 620 -203
rect 655 -208 661 -137
rect 684 -181 689 -99
rect 735 -114 739 -99
rect 692 -121 716 -114
rect 770 -117 774 -99
rect 801 -110 858 -103
rect 807 -116 811 -110
rect 840 -116 844 -110
rect 698 -127 702 -121
rect 706 -181 710 -167
rect 684 -185 699 -181
rect 706 -185 721 -181
rect 706 -189 710 -185
rect 616 -211 661 -208
rect 716 -195 721 -185
rect 731 -182 735 -161
rect 782 -157 800 -153
rect 739 -170 743 -161
rect 796 -170 800 -157
rect 815 -170 819 -156
rect 848 -170 852 -156
rect 739 -174 808 -170
rect 815 -174 841 -170
rect 848 -174 860 -170
rect 771 -182 775 -174
rect 731 -186 739 -182
rect 751 -195 755 -190
rect 716 -199 755 -195
rect 616 -212 669 -211
rect 612 -223 616 -219
rect 648 -223 652 -212
rect 658 -216 669 -212
rect 698 -218 702 -209
rect 798 -193 802 -174
rect 815 -178 819 -174
rect 848 -178 852 -174
rect 795 -196 802 -193
rect 783 -218 787 -210
rect 807 -218 811 -198
rect 840 -218 844 -198
rect 561 -227 576 -223
rect 583 -227 616 -223
rect 692 -226 859 -218
rect 583 -231 587 -227
rect 470 -240 518 -237
rect 273 -251 277 -245
rect 306 -251 310 -245
rect 259 -258 316 -251
rect 343 -262 347 -244
rect 401 -247 425 -240
rect 428 -246 518 -240
rect 378 -262 382 -247
rect 428 -262 433 -246
rect 470 -249 518 -246
rect 343 -266 433 -262
rect 470 -265 518 -252
rect 575 -260 579 -251
rect 644 -260 648 -231
rect 569 -268 669 -260
rect 258 -277 425 -269
rect 648 -275 661 -271
rect 273 -297 277 -277
rect 306 -297 310 -277
rect 330 -285 334 -277
rect 315 -302 322 -299
rect 265 -321 269 -317
rect 298 -321 302 -317
rect 315 -321 319 -302
rect 415 -286 419 -277
rect 362 -300 401 -296
rect 362 -305 366 -300
rect 378 -313 386 -309
rect 342 -321 346 -313
rect 257 -325 269 -321
rect 276 -325 302 -321
rect 309 -325 378 -321
rect 265 -339 269 -325
rect 298 -339 302 -325
rect 317 -338 321 -325
rect 374 -334 378 -325
rect 317 -342 335 -338
rect 382 -334 386 -313
rect 396 -310 401 -300
rect 561 -279 621 -275
rect 407 -310 411 -306
rect 396 -314 411 -310
rect 418 -314 433 -310
rect 407 -328 411 -314
rect 415 -374 419 -368
rect 273 -385 277 -379
rect 306 -385 310 -379
rect 259 -392 316 -385
rect 343 -396 347 -378
rect 401 -381 425 -374
rect 378 -396 382 -381
rect 428 -382 433 -314
rect 561 -361 566 -279
rect 644 -292 648 -283
rect 569 -301 593 -294
rect 602 -295 648 -292
rect 608 -301 612 -295
rect 575 -307 579 -301
rect 583 -361 587 -347
rect 616 -346 620 -341
rect 655 -346 661 -275
rect 616 -349 661 -346
rect 616 -350 670 -349
rect 612 -361 616 -357
rect 648 -361 652 -350
rect 658 -354 670 -350
rect 561 -365 576 -361
rect 583 -365 616 -361
rect 583 -369 587 -365
rect 470 -382 518 -377
rect 428 -388 518 -382
rect 428 -396 433 -388
rect 470 -390 518 -388
rect 343 -400 433 -396
rect 470 -406 518 -393
rect 575 -398 579 -389
rect 644 -398 648 -369
rect 569 -406 670 -398
<< metal2 >>
rect 208 655 302 662
rect 208 651 216 655
rect 693 654 722 659
rect 726 654 755 659
rect 759 654 788 659
rect 792 654 821 659
rect 825 654 842 659
rect 838 650 842 654
rect 523 625 552 630
rect 556 625 585 630
rect 589 625 618 630
rect 622 625 639 630
rect 635 621 639 625
rect 386 604 415 609
rect 419 604 448 609
rect 452 604 469 609
rect 465 600 469 604
rect 220 517 314 524
rect 220 513 228 517
rect 402 462 431 467
rect 435 462 464 467
rect 468 462 485 467
rect 539 464 568 469
rect 572 464 601 469
rect 605 464 634 469
rect 638 464 655 469
rect 481 458 485 462
rect 651 460 655 464
rect 715 409 719 458
rect 715 405 740 409
rect 698 394 715 398
rect 719 394 744 398
rect 748 394 777 398
rect 781 394 787 398
rect 273 379 367 386
rect 867 381 871 430
rect 273 375 281 379
rect 867 377 892 381
rect 337 368 577 373
rect 458 301 487 306
rect 491 301 520 306
rect 524 301 541 306
rect 537 297 541 301
rect 273 241 367 248
rect 273 237 281 241
rect 572 165 576 368
rect 830 366 846 370
rect 850 366 867 370
rect 871 366 896 370
rect 900 366 929 370
rect 933 366 939 370
rect 740 333 834 340
rect 740 329 748 333
rect 601 270 605 319
rect 806 271 812 278
rect 601 266 626 270
rect 768 265 825 271
rect 819 260 825 265
rect 605 255 630 259
rect 634 255 663 259
rect 667 255 673 259
rect 703 170 797 177
rect 703 166 711 170
rect 488 160 679 165
rect 488 133 492 160
rect 462 117 491 121
rect 495 117 501 121
rect 324 85 330 90
rect 324 79 381 85
rect 385 79 463 85
rect 337 72 343 79
rect 455 21 463 79
rect 633 21 638 114
rect 673 72 679 160
rect 769 108 775 115
rect 731 102 788 108
rect 782 97 788 102
rect 669 64 679 72
rect 401 17 409 21
rect 315 10 409 17
rect 455 14 507 21
rect 515 16 638 21
rect 702 24 796 31
rect 702 20 710 24
rect 324 -49 330 -44
rect 324 -55 381 -49
rect 385 -55 452 -49
rect 337 -62 343 -55
rect 401 -117 409 -113
rect 315 -124 409 -117
rect 443 -116 452 -55
rect 628 -116 635 -23
rect 768 -38 774 -31
rect 730 -44 787 -38
rect 781 -49 787 -44
rect 707 -110 801 -103
rect 707 -114 715 -110
rect 443 -123 504 -116
rect 514 -121 635 -116
rect 325 -183 331 -178
rect 325 -189 382 -183
rect 386 -189 451 -183
rect 338 -196 344 -189
rect 402 -251 410 -247
rect 316 -258 410 -251
rect 444 -254 451 -189
rect 637 -254 642 -161
rect 773 -172 779 -165
rect 735 -178 792 -172
rect 786 -183 792 -178
rect 444 -259 509 -254
rect 516 -259 642 -254
rect 325 -317 331 -312
rect 325 -323 382 -317
rect 386 -323 450 -317
rect 338 -330 344 -323
rect 402 -385 410 -381
rect 316 -392 410 -385
rect 442 -394 450 -323
rect 635 -393 640 -299
rect 442 -400 509 -394
rect 516 -397 640 -393
<< metal3 >>
rect 502 47 572 55
rect 502 32 509 47
rect 506 -88 571 -83
rect 506 -102 513 -88
rect 510 -229 574 -223
rect 510 -240 515 -229
rect 507 -367 575 -361
rect 507 -379 514 -367
<< pad >>
rect 302 655 310 662
rect 689 654 694 659
rect 722 654 727 659
rect 755 654 760 659
rect 788 654 793 659
rect 821 654 826 659
rect 208 644 216 651
rect 838 646 843 651
rect 519 625 524 630
rect 552 625 557 630
rect 585 625 590 630
rect 618 625 623 630
rect 635 617 640 622
rect 382 604 387 609
rect 415 604 420 609
rect 448 604 453 609
rect 465 596 470 601
rect 314 517 322 524
rect 220 506 228 513
rect 398 462 403 467
rect 431 462 436 467
rect 464 462 469 467
rect 535 464 540 469
rect 568 464 573 469
rect 601 464 606 469
rect 634 464 639 469
rect 481 454 486 459
rect 651 456 656 461
rect 719 454 724 459
rect 871 426 876 431
rect 740 405 745 410
rect 694 394 699 399
rect 715 394 720 399
rect 744 394 749 399
rect 777 394 782 399
rect 787 394 792 399
rect 367 379 375 386
rect 892 377 897 382
rect 273 368 281 375
rect 330 368 337 375
rect 826 366 831 371
rect 846 366 851 371
rect 867 366 872 371
rect 896 366 901 371
rect 929 366 934 371
rect 939 366 944 371
rect 834 333 842 340
rect 740 322 748 329
rect 605 315 610 320
rect 454 301 459 306
rect 487 301 492 306
rect 520 301 525 306
rect 537 293 542 298
rect 626 266 631 271
rect 764 265 769 271
rect 601 255 606 260
rect 630 255 635 260
rect 663 255 668 260
rect 673 255 678 260
rect 367 241 375 248
rect 273 230 281 237
rect 797 170 805 177
rect 703 159 711 166
rect 488 130 493 135
rect 458 117 463 122
rect 491 117 496 122
rect 501 117 506 122
rect 633 114 641 122
rect 727 102 732 108
rect 381 79 386 85
rect 661 64 669 72
rect 572 47 580 55
rect 502 30 510 38
rect 401 21 409 28
rect 796 24 804 31
rect 307 10 315 17
rect 507 14 515 22
rect 702 13 710 20
rect 628 -23 635 -16
rect 726 -44 731 -38
rect 381 -55 386 -49
rect 570 -90 577 -83
rect 401 -113 409 -106
rect 504 -108 514 -99
rect 801 -110 809 -103
rect 307 -124 315 -117
rect 504 -124 514 -115
rect 707 -121 715 -114
rect 637 -161 644 -154
rect 731 -178 736 -172
rect 382 -189 387 -183
rect 573 -229 580 -222
rect 402 -247 410 -240
rect 508 -244 515 -237
rect 308 -258 316 -251
rect 509 -259 516 -252
rect 635 -299 642 -292
rect 382 -323 387 -317
rect 573 -367 580 -360
rect 402 -381 410 -374
rect 507 -384 514 -377
rect 308 -392 316 -385
rect 509 -400 516 -393
<< labels >>
rlabel metal1 580 -299 580 -299 5 vdd
rlabel metal1 575 -402 575 -402 1 gnd
rlabel metal1 580 -161 580 -161 5 vdd
rlabel metal1 575 -264 575 -264 1 gnd
rlabel metal1 577 -23 577 -23 5 vdd
rlabel metal1 572 -126 572 -126 1 gnd
rlabel metal1 484 32 484 32 1 a0
rlabel metal1 485 15 485 15 1 b0
rlabel metal1 492 -103 492 -103 1 a1
rlabel metal1 493 -243 493 -243 1 a2
rlabel metal1 497 -383 497 -383 1 a3
rlabel metal1 493 -399 493 -399 1 b3
rlabel metal1 496 -257 496 -257 1 b2
rlabel metal1 488 -121 488 -121 1 b1
rlabel metal1 637 14 637 14 1 gnd
rlabel metal1 580 115 580 115 5 vdd
rlabel metal1 418 129 418 129 5 gnd
rlabel metal1 304 15 304 15 1 vdd
rlabel metal1 413 26 413 26 1 vdd
rlabel metal1 261 79 261 79 3 p0
rlabel metal1 261 -55 261 -55 1 p1
rlabel metal1 413 -108 413 -108 1 vdd
rlabel metal1 304 -119 304 -119 1 vdd
rlabel metal1 418 -5 418 -5 5 gnd
rlabel metal1 419 -139 419 -139 5 gnd
rlabel metal1 305 -253 305 -253 1 vdd
rlabel metal1 414 -242 414 -242 1 vdd
rlabel metal1 259 -188 259 -188 1 p2
rlabel metal1 419 -273 419 -273 5 gnd
rlabel metal1 305 -387 305 -387 1 vdd
rlabel metal1 414 -376 414 -376 1 vdd
rlabel metal1 261 -322 261 -322 1 p3
rlabel metal1 411 243 411 243 5 vdd
rlabel metal1 378 243 378 243 5 vdd
rlabel metal1 269 232 269 232 5 vdd
rlabel metal1 332 237 332 237 1 cin
rlabel metal1 422 178 422 178 1 pocin
rlabel metal1 517 193 517 193 5 vdd
rlabel metal1 511 98 511 98 1 gnd
rlabel metal1 530 127 530 127 1 c1
rlabel metal1 418 267 418 267 5 gnd
rlabel metal1 411 381 411 381 5 vdd
rlabel metal1 378 381 378 381 5 vdd
rlabel metal1 269 370 269 370 5 vdd
rlabel metal1 424 317 424 317 1 p1g0
rlabel metal1 545 227 545 227 1 gnd
rlabel metal1 507 363 507 363 5 vdd
rlabel metal1 451 292 451 292 1 p1
rlabel metal1 475 292 475 292 1 p0
rlabel metal1 489 285 489 285 1 cin
rlabel metal1 216 508 216 508 5 vdd
rlabel metal1 325 519 325 519 5 vdd
rlabel metal1 358 519 358 519 5 vdd
rlabel metal1 211 405 211 405 1 gnd
rlabel metal1 451 524 451 524 5 vdd
rlabel metal1 489 388 489 388 1 gnd
rlabel metal1 659 390 659 390 1 gnd
rlabel metal1 621 526 621 526 5 vdd
rlabel metal1 797 375 797 375 1 gnd
rlabel metal1 803 470 803 470 5 vdd
rlabel metal1 533 443 533 443 1 p2
rlabel metal1 565 446 565 446 1 p1
rlabel metal1 589 447 589 447 1 p0
rlabel metal1 602 442 602 442 1 cin
rlabel metal1 680 458 680 458 1 p2p1p0c0
rlabel metal1 691 407 691 407 1 g2
rlabel metal1 713 408 713 408 1 p2g1g0
rlabel pad 742 408 742 408 1 p2p1p0c0
rlabel metal1 202 444 202 444 3 p2
rlabel metal1 269 514 269 514 1 g1
rlabel metal1 368 454 368 454 1 p2g1
rlabel metal1 396 449 396 449 1 p2
rlabel metal1 418 449 418 449 1 p1
rlabel metal1 434 441 434 441 1 g0
rlabel metal1 511 457 511 457 1 p2p1g0
rlabel metal1 775 409 775 409 1 p2g1
rlabel metal1 815 404 815 404 7 c3
rlabel metal1 204 646 204 646 5 vdd
rlabel metal1 346 657 346 657 5 vdd
rlabel metal1 199 543 199 543 1 gnd
rlabel metal1 435 666 435 666 5 vdd
rlabel metal1 473 530 473 530 1 gnd
rlabel metal1 605 687 605 687 5 vdd
rlabel metal1 643 551 643 551 1 gnd
rlabel metal1 808 716 808 716 5 vdd
rlabel metal1 846 580 846 580 1 gnd
rlabel metal1 949 347 949 347 1 gnd
rlabel metal1 955 442 955 442 5 vdd
rlabel metal1 192 583 192 583 1 p3
rlabel metal1 264 652 264 652 1 g2
rlabel metal1 359 593 359 593 1 p3g2
rlabel metal1 379 591 379 591 1 p3
rlabel metal1 402 591 402 591 1 p2
rlabel metal1 418 585 418 585 1 g1
rlabel metal1 494 597 494 597 1 p3p2g1
rlabel metal1 516 599 516 599 1 p3
rlabel metal1 550 603 550 603 1 p2
rlabel metal1 586 604 586 604 1 g0
rlabel metal1 666 619 666 619 1 p3p2p1g0
rlabel metal1 686 633 686 633 1 p3
rlabel metal1 720 624 720 624 1 p2
rlabel metal1 753 631 753 631 1 p1
rlabel metal1 775 638 775 638 1 p0
rlabel metal1 790 636 790 636 1 cin
rlabel metal1 867 648 867 648 1 p3p2p1p0c0
rlabel metal1 824 398 824 398 1 g3
rlabel metal1 843 395 843 395 1 p3g2
rlabel metal1 864 395 864 395 1 p3p2g1
rlabel metal1 928 379 928 379 1 p3p2p1p0c0
rlabel metal1 966 376 966 376 7 c4
rlabel metal1 736 324 736 324 5 vdd
rlabel metal1 845 335 845 335 5 vdd
rlabel metal1 878 335 878 335 5 vdd
rlabel metal1 731 221 731 221 1 gnd
rlabel metal1 726 260 726 260 1 p0
rlabel pad 766 268 766 268 1 cin
rlabel metal1 892 271 892 271 1 s0
rlabel pad 894 380 894 380 1 p3p2p1g0
rlabel metal1 570 295 570 295 1 p1p0c0
rlabel pad 489 131 489 131 1 g0
rlabel metal1 683 236 683 236 1 gnd
rlabel metal1 689 331 689 331 5 vdd
rlabel metal1 698 265 698 265 1 c2
rlabel metal1 598 272 598 272 1 g1
rlabel pad 628 267 628 267 1 p1g0
rlabel metal1 661 268 661 268 1 p1p0c0
rlabel metal1 573 612 573 612 1 p1
rlabel metal1 655 -72 655 -72 1 g1
rlabel metal1 663 -213 663 -213 1 g2
rlabel metal1 666 -351 666 -351 1 g3
rlabel metal1 699 161 699 161 5 vdd
rlabel metal1 808 172 808 172 5 vdd
rlabel metal1 841 172 841 172 5 vdd
rlabel metal1 694 58 694 58 1 gnd
rlabel metal1 852 108 852 108 1 s1
rlabel metal1 686 97 686 97 1 p1
rlabel pad 728 105 728 105 1 c1
rlabel metal1 698 15 698 15 5 vdd
rlabel metal1 807 26 807 26 5 vdd
rlabel metal1 840 26 840 26 5 vdd
rlabel metal1 693 -88 693 -88 1 gnd
rlabel metal1 852 -38 852 -38 1 s2
rlabel metal1 682 -49 682 -49 1 p2
rlabel pad 728 -41 728 -41 1 c2
rlabel metal1 698 -222 698 -222 1 gnd
rlabel metal1 845 -108 845 -108 5 vdd
rlabel metal1 812 -108 812 -108 5 vdd
rlabel metal1 703 -119 703 -119 5 vdd
rlabel metal1 855 -171 855 -171 7 s3
rlabel metal1 688 -184 688 -184 1 p3
rlabel pad 733 -176 733 -176 1 c3
rlabel metal2 672 67 672 67 1 g0
rlabel metal1 658 68 658 68 1 g0
<< end >>
