magic
tech scmos
timestamp 1731796585
<< nwell >>
rect -216 -43 -160 -18
rect -147 -43 -91 -18
rect -85 -43 -29 -18
rect -216 -73 -160 -49
rect -23 -70 7 -14
<< ntransistor >>
rect -118 -56 -98 -54
rect -56 -56 -36 -54
rect -214 -87 -194 -85
rect -144 -87 -124 -85
rect -82 -87 -62 -85
rect -6 -110 -4 -90
<< ptransistor >>
rect -206 -31 -166 -29
rect -137 -31 -97 -29
rect -75 -31 -35 -29
rect -206 -62 -166 -60
rect -6 -60 -4 -20
<< ndiffusion >>
rect -118 -54 -98 -53
rect -118 -57 -98 -56
rect -56 -54 -36 -53
rect -56 -57 -36 -56
rect -214 -85 -194 -84
rect -214 -88 -194 -87
rect -144 -85 -124 -84
rect -82 -85 -62 -84
rect -144 -88 -124 -87
rect -82 -88 -62 -87
rect -7 -110 -6 -90
rect -4 -110 -3 -90
<< pdiffusion >>
rect -206 -29 -166 -28
rect -206 -32 -166 -31
rect -137 -29 -97 -28
rect -137 -32 -97 -31
rect -75 -29 -35 -28
rect -75 -32 -35 -31
rect -206 -60 -166 -59
rect -7 -60 -6 -20
rect -4 -60 -3 -20
rect -206 -63 -166 -62
<< ndcontact >>
rect -118 -53 -98 -49
rect -56 -53 -36 -49
rect -118 -61 -98 -57
rect -56 -61 -36 -57
rect -214 -84 -194 -80
rect -144 -84 -124 -80
rect -82 -84 -62 -80
rect -214 -92 -194 -88
rect -144 -92 -124 -88
rect -82 -92 -62 -88
rect -11 -110 -7 -90
rect -3 -110 1 -90
<< pdcontact >>
rect -206 -28 -166 -24
rect -137 -28 -97 -24
rect -75 -28 -35 -24
rect -206 -36 -166 -32
rect -137 -36 -97 -32
rect -75 -36 -35 -32
rect -206 -59 -166 -55
rect -11 -60 -7 -20
rect -3 -60 1 -20
rect -206 -67 -166 -63
<< polysilicon >>
rect -6 -20 -4 -17
rect -216 -31 -206 -29
rect -166 -31 -163 -29
rect -147 -31 -137 -29
rect -97 -31 -94 -29
rect -84 -31 -75 -29
rect -35 -31 -32 -29
rect -121 -56 -118 -54
rect -98 -56 -95 -54
rect -59 -56 -56 -54
rect -36 -56 -33 -54
rect -216 -62 -206 -60
rect -166 -62 -163 -60
rect -217 -87 -214 -85
rect -194 -87 -191 -85
rect -147 -87 -144 -85
rect -124 -87 -121 -85
rect -85 -87 -82 -85
rect -62 -87 -59 -85
rect -6 -90 -4 -60
rect -6 -113 -4 -110
<< polycontact >>
rect -220 -32 -216 -28
rect -151 -32 -147 -28
rect -88 -32 -84 -28
rect -125 -57 -121 -53
rect -63 -57 -59 -53
rect -220 -63 -216 -59
rect -221 -88 -217 -84
rect -151 -88 -147 -84
rect -89 -87 -85 -83
rect -10 -86 -6 -82
<< metal1 >>
rect -160 -14 7 -11
rect -160 -24 -157 -14
rect -100 -24 -97 -14
rect -40 -24 -37 -14
rect -11 -20 -7 -14
rect -166 -28 -157 -24
rect -236 -32 -220 -28
rect -152 -32 -151 -28
rect -236 -84 -233 -32
rect -169 -55 -166 -36
rect -101 -43 -98 -36
rect -88 -43 -85 -32
rect -101 -46 -85 -43
rect -39 -43 -36 -36
rect -39 -46 -25 -43
rect -101 -49 -98 -46
rect -160 -56 -125 -53
rect -229 -63 -220 -59
rect -213 -67 -206 -63
rect -213 -71 -210 -67
rect -160 -71 -157 -56
rect -213 -74 -157 -71
rect -101 -73 -98 -61
rect -213 -80 -210 -74
rect -144 -76 -98 -73
rect -144 -80 -141 -76
rect -90 -83 -87 -46
rect -39 -49 -36 -46
rect -71 -56 -63 -53
rect -39 -73 -36 -61
rect -82 -76 -36 -73
rect -82 -80 -79 -76
rect -236 -88 -221 -84
rect -152 -88 -151 -84
rect -90 -87 -89 -83
rect -29 -82 -25 -46
rect -3 -82 1 -60
rect -29 -86 -10 -82
rect -3 -86 7 -82
rect -194 -92 -181 -88
rect -124 -92 -111 -88
rect -62 -92 -49 -88
rect -3 -90 1 -86
rect -184 -95 -181 -92
rect -114 -95 -111 -92
rect -52 -95 -49 -92
rect -34 -95 -23 -94
rect -184 -98 -23 -95
rect -27 -119 -23 -98
rect -11 -119 -7 -110
rect -27 -122 7 -119
<< metal2 >>
rect -155 -58 -150 -29
rect -224 -60 -150 -58
rect -68 -60 -65 -53
rect -224 -63 -63 -60
rect -155 -64 -63 -63
rect -155 -84 -150 -64
<< pad >>
rect -155 -35 -150 -29
rect -71 -57 -65 -52
rect -224 -63 -219 -58
rect -155 -88 -150 -82
<< labels >>
rlabel metal1 -235 -51 -235 -51 3 d
rlabel metal1 -184 -91 -184 -91 7 gnd
rlabel metal1 -114 -91 -114 -91 7 gnd
rlabel metal1 -226 -61 -226 -61 3 clk
rlabel metal1 -52 -91 -52 -91 7 gnd
rlabel metal1 -6 -12 -6 -12 5 vdd
rlabel metal1 -10 -120 -10 -120 1 gnd
rlabel metal1 1 -84 1 -84 1 q
rlabel metal1 -18 -83 -18 -83 1 qbar
<< end >>
