* SPICE3 file created from or4.ext - technology: scmos

.option scale=1u

M1000 vdd d a_n75_82# w_n80_103# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1001 ybar b gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 ybar a gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 ybar d gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1004 ybar c gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 ybar c a_n75_7# w_n81_1# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 y ybar vdd w_n16_0# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 a_n75_47# b a_n75_7# w_n81_34# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 a_n75_82# a a_n75_47# w_n81_69# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1009 y ybar gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
C0 ybar w_n16_0# 1.014f
C1 a_n75_7# w_n81_1# 2.444f
C2 w_n80_103# a_n75_82# 1.41f
C3 w_n16_0# vdd 1.128f
C4 a_n75_47# w_n81_34# 1.41f
C5 w_n16_0# y 1.88f
C6 a_n75_7# w_n81_34# 1.128f
C7 w_n80_103# d 1.482f
C8 w_n81_69# a_n75_47# 1.41f
C9 ybar gnd 2.424f
C10 c w_n81_1# 2.312f
C11 w_n81_69# a_n75_82# 1.598f
C12 ybar w_n81_1# 1.88f
C13 b w_n81_34# 1.482f
C14 w_n80_103# vdd 1.88f
C15 w_n81_69# a 1.482f
C16 gnd 0 19.834f **FLOATING
C17 y 0 4.324f **FLOATING
C18 c 0 8.299999f **FLOATING
C19 a_n75_7# 0 4.888f **FLOATING
C20 b 0 14.034f **FLOATING
C21 ybar 0 22.275f **FLOATING
C22 a_n75_47# 0 2.585f **FLOATING
C23 a 0 25.962f **FLOATING
C24 a_n75_82# 0 2.35f **FLOATING
C25 d 0 36.49f **FLOATING
C26 vdd 0 23.03f **FLOATING
