* SPICE3 file created from testing_withoutbuffer.ext - technology: scmos

.option scale=90n

M1000 a_594_537# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1001 a_582_n389# a3 vdd w_569_n357# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1002 a_239_604# p3 g2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 gnd a_325_n314# a_303_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1004 gnd a_303_n382# a_270_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 a_218_418# p2 vdd w_205_450# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 a_825_350# g3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1007 a_617_285# p1p0c0 a_617_278# w_611_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 c1 a_445_147# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1009 p3p2p1g0 a_518_635# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1010 a_731_424# p2g1 a_731_417# w_725_411# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1011 a_662_239# p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 gnd a_270_n248# p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 gnd a_269_20# p0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 a_594_556# p2 a_594_537# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 g3 a_582_n389# b3 w_602_n351# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1016 g2 a_582_n251# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1017 a_490_101# g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1018 s1 a_810_82# vdd w_830_114# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_594_575# p1 a_594_556# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1020 p2g1 a_327_429# vdd w_347_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1021 a_440_412# p1 a_440_393# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 p1p0c0 a_453_311# vdd w_544_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a3 a_338_n335# a_303_n382# w_329_n384# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1024 s2 a_809_n64# vdd w_829_n32# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1025 a_518_635# p3 vdd w_505_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1026 a_731_457# a_724_454# a_731_417# w_725_444# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1027 b2 a2 a_303_n248# w_368_n246# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1028 gnd a_303_n248# a_270_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1029 p3p2g1 a_381_614# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 p2p1p0c0 a_534_474# vdd w_658_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 a_610_395# p1 a_610_377# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1032 gnd a_325_n180# a_303_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1033 a_518_635# g0 a_594_575# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1034 a_705_n209# p3 vdd w_692_n177# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 vdd a0 a_345_92# w_400_28# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1036 vdd a_302_20# a_269_20# w_291_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1037 s3 a_814_n198# vdd w_834_n166# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1038 a_346_n176# b2 a_303_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1039 a_734_119# c1 a_701_71# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1040 a_866_350# p3p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1041 a_847_245# a_771_282# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 a_304_190# a_271_142# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1043 a_884_498# p3g2 a_883_464# w_878_485# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1044 a_733_n27# c2 a_700_n75# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1045 a_731_492# p2g1g0 a_731_457# w_725_479# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 g3 a3 b3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1047 a_315_567# a_239_604# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 a_582_n251# a2 vdd w_569_n219# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 p3g2 a_315_567# vdd w_335_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 vdd g3 a_884_498# w_879_518# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1051 a_895_350# a_892_373# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1052 pocin a_380_153# vdd w_400_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 vdd a_269_20# p0 w_258_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1054 a_218_418# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1055 a_380_153# a_304_190# vdd w_367_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 b1 a1 a_302_n114# w_367_n112# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 a_928_350# p3p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1058 a_271_280# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 a_814_n198# a_738_n161# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 p3p2p1g0 a_518_635# vdd w_642_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_239_604# a_206_556# g2 w_226_594# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_304_190# a_271_142# cin w_291_180# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 g2 a_582_n251# b2 w_602_n213# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1064 g1 a_579_n113# b1 w_599_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1065 a_582_25# a0 vdd w_569_57# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1066 a_734_119# a_769_115# p1 w_760_117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1067 c3 a_731_424# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1068 p2p1g0 a_397_472# vdd w_488_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_440_393# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 g1 a_579_n113# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1071 a_688_664# p0 vdd w_774_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1072 a_457_101# pocin gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 p2g1 a_327_429# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_629_239# a_626_262# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1075 a_327_429# a_251_466# vdd w_314_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1076 a_700_n75# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1077 a_688_664# cin vdd w_807_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1078 a_776_378# p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1079 a_251_466# p2 g1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1080 a_705_n209# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1081 a_346_n310# b3 a_303_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1082 a_810_82# a_734_119# vdd w_797_114# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1083 a_738_234# p0 vdd w_725_266# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1084 p3p2g1 a_381_614# vdd w_472_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1085 a_809_n64# a_733_n27# vdd w_796_n32# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_206_556# p3 vdd w_193_588# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1087 a_424_535# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1088 s1 a_810_82# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1089 a_610_377# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 s0 a_847_245# vdd w_867_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_582_n389# a3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 vdd a2 a_346_n176# w_401_n240# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 g2 a2 b2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1094 c4 a_883_396# vdd w_942_382# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 a_738_n161# p3 c3 w_725_n171# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1096 a_810_82# a_734_119# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1097 a_424_554# p2 a_424_535# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_453_311# p0 vdd w_473_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1099 a_315_567# a_239_604# vdd w_302_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 p3p2p1p0c0 a_688_664# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1101 a_771_282# p0 cin w_758_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1102 a_271_142# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1103 g1 a1 b1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1104 a_534_474# cin vdd w_620_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_534_474# p0 vdd w_587_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_453_311# cin vdd w_506_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1107 a_271_280# p1 vdd w_258_312# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_381_614# g1 a_424_554# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 a_883_429# a_876_426# a_883_389# w_877_416# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1110 a_714_378# p2g1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 a_701_71# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 c1 a_445_147# vdd w_504_133# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1113 a_304_328# a_271_280# g0 w_291_318# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 a_845_350# p3g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1115 a_688_664# p1 vdd w_741_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1116 a_797_604# p0 a_797_585# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1117 vdd a_269_n114# p1 w_258_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1118 p1g0 a_380_291# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 s2 a_809_n64# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1120 a_345_n42# b1 a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1121 a_327_429# a_251_466# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1122 a_733_n27# p2 c2 w_720_n37# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 a_743_378# a_740_401# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1124 a_380_291# a_304_328# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 c2 a_617_285# vdd w_676_271# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1126 b3 a3 a_303_n382# w_368_n380# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1127 a1 a_337_n67# a_302_n114# w_328_n116# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1128 gnd a_324_n46# a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1129 gnd a_324_88# a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1130 vdd a3 a_346_n310# w_401_n374# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1131 g0 a_582_25# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1132 p1p0c0 a_453_311# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_345_92# b0 a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1134 a_688_664# cin a_797_604# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1135 vdd g2 a_731_492# w_726_513# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1136 a_883_464# p3p2g1 a_883_429# w_877_451# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1137 a_693_378# g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1138 s3 a_814_n198# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1139 a_304_328# p1 g0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1140 a_771_282# a_819_257# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1141 a_518_635# p1 vdd w_571_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_397_472# g0 vdd w_450_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_579_n113# a1 vdd w_566_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 a_797_547# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1145 a_496_251# p0 a_496_232# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_518_635# g0 vdd w_604_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1147 a_883_396# p3p2p1p0c0 a_883_389# w_877_383# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1148 p2p1p0c0 a_534_474# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1149 a_847_245# a_771_282# vdd w_834_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1150 vdd a_270_n248# p2 w_259_n251# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 a_579_n113# a1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1152 a_239_604# a_206_556# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1153 a_797_566# p2 a_797_547# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1154 a_453_311# cin a_496_251# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 a_453_311# p1 vdd w_440_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 gnd a3 a_346_n310# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_534_474# p1 vdd w_554_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1158 a_304_328# a_271_280# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1159 a_445_147# g0 a_445_140# w_439_134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1160 a_797_585# p1 a_797_566# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 a_733_n27# a_781_n52# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 gnd a_302_n114# a_269_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1163 gnd a_269_n114# p1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 vdd a_303_n248# a_270_n248# w_292_n251# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1165 a_381_614# g1 vdd w_434_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1166 pocin a_380_153# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1167 a_380_153# a_304_190# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1168 a_688_664# p3 vdd w_675_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1169 p1g0 a_380_291# vdd w_400_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1170 c2 a_617_285# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 a0 a_337_67# a_302_20# w_328_18# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1172 g0 a0 b0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1173 a_380_291# a_304_328# vdd w_367_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 vdd a_270_n382# p3 w_259_n385# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1175 a_582_25# a0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1176 a_701_71# p1 vdd w_688_103# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1177 a_688_664# p2 vdd w_708_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1178 p2p1g0 a_397_472# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1179 gnd a2 a_346_n176# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1180 vdd pocin a_445_140# w_439_167# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1181 a_809_n64# a_733_n27# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1182 c3 a_731_424# vdd w_790_410# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 a_304_190# p0 cin Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1184 a_734_119# p1 c1 w_721_109# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1185 a_251_466# a_218_418# g1 w_238_456# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 vdd a1 a_345_n42# w_400_n106# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1187 a_814_n198# a_738_n161# vdd w_801_n166# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1188 a_397_472# g0 a_440_412# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 a_738_n161# c3 a_705_n209# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1190 g3 a_582_n389# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1191 a_738_n161# a_773_n165# p3 w_764_n163# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1192 a_397_472# p2 vdd w_384_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1193 vdd a_302_n114# a_269_n114# w_291_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 a_617_318# a_610_315# a_617_278# w_611_305# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1195 a_771_282# a_806_278# p0 w_797_280# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_738_234# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1197 vdd a_303_n382# a_270_n382# w_292_n385# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_518_635# p2 vdd w_538_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1199 a_496_232# p1 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 b0 a0 a_302_20# w_367_22# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1201 a_397_472# p1 vdd w_417_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 a_700_n75# p2 vdd w_687_n43# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_734_119# a_782_94# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1204 a_206_556# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1205 gnd a_270_n382# p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 p3p2p1p0c0 a_688_664# vdd w_845_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 a_610_414# p0 a_610_395# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1208 a_582_n251# a2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1209 a_534_474# p2 vdd w_521_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1210 a_271_142# p0 vdd w_258_174# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1211 s0 a_847_245# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1212 vdd g1 a_617_318# w_611_340# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 c4 a_883_396# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 gnd a1 a_345_n42# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1215 gnd a0 a_345_92# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 gnd a_302_20# a_269_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1217 a_381_614# p2 vdd w_401_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1218 a2 a_338_n201# a_303_n248# w_329_n250# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1219 a_733_n27# a_768_n31# p2 w_759_n29# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1220 a_251_466# a_218_418# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1221 a_534_474# cin a_610_414# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1222 a_771_282# cin a_738_234# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1223 a_381_614# p3 vdd w_368_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1224 p3g2 a_315_567# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1225 a_600_239# g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1226 a_738_n161# a_786_n186# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1227 g0 a_582_25# b0 w_602_63# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 a_809_n64# vdd 0.441416f
C1 a_733_n27# gnd 0.396612f
C2 b2 a_303_n248# 0.599413f
C3 w_521_464# p2 0.026794f
C4 w_675_654# p3 0.026794f
C5 a_617_285# c2 0.060798f
C6 a_731_417# p2p1p0c0 0.004158f
C7 w_292_n251# a_270_n248# 0.013216f
C8 w_368_n246# b2 0.014021f
C9 w_401_n240# a2 0.028034f
C10 w_569_57# vdd 0.008451f
C11 a_700_n75# p2 0.060798f
C12 a_251_466# a_218_418# 0.003752f
C13 w_439_134# pocin 1.21e-19
C14 a_490_101# gnd 0.247451f
C15 a_582_25# vdd 0.439883f
C16 w_205_450# p2 0.028034f
C17 w_571_625# a_518_635# 0.028268f
C18 a_610_377# p2 0.013746f
C19 a_883_396# g3 1.39e-20
C20 p1 a_734_119# 0.413834f
C21 w_439_167# vdd 0.010186f
C22 a_810_82# gnd 0.248155f
C23 a0 vdd 0.228122f
C24 w_877_451# p3p2g1 0.036563f
C25 w_845_654# p3p2p1p0c0 0.013216f
C26 w_725_444# a_731_417# 0.008113f
C27 a_731_492# vdd 0.41238f
C28 w_450_462# g0 0.026794f
C29 w_758_272# vdd 6.13e-19
C30 a_797_585# p1 0.013746f
C31 w_611_305# p1g0 2.18e-19
C32 a_883_396# a_845_350# 0.002189f
C33 a_380_153# gnd 0.248155f
C34 a_271_142# vdd 0.439891f
C35 w_797_280# cin 1.23e-19
C36 w_291_180# a_304_190# 0.019526f
C37 w_867_277# s0 0.013216f
C38 w_725_479# p2g1g0 0.036563f
C39 w_878_485# a_883_464# 0.009864f
C40 a_594_537# p3 0.013746f
C41 a_346_n310# gnd 0.20619f
C42 a_582_n389# vdd 0.439883f
C43 a_304_328# g0 0.753587f
C44 w_473_301# vdd 0.008451f
C45 w_796_n32# a_809_n64# 0.013216f
C46 b1 a_302_n114# 0.599413f
C47 s0 gnd 0.20619f
C48 a_626_262# p1g0 2.36e-20
C49 a_768_n31# c2 5.8e-19
C50 a_733_n27# a_700_n75# 0.20619f
C51 w_506_301# cin 0.026794f
C52 a1 a_345_n42# 0.060798f
C53 g1 a_579_n113# 0.003752f
C54 p0 vdd 0.678634f
C55 a_688_664# gnd 0.042086f
C56 p0 a_496_232# 0.013746f
C57 w_658_464# a_534_474# 0.027163f
C58 w_725_479# a_731_492# 0.01128f
C59 a_397_472# p2 0.002443f
C60 a_518_635# vdd 1.76176f
C61 w_878_485# a_884_498# 0.01128f
C62 a_206_556# p3 0.060798f
C63 b3 a_582_n389# 0.00288f
C64 a3 a_338_n335# 0.014473f
C65 a_731_424# a_776_378# 0.029681f
C66 g3 vdd 0.002989f
C67 a_786_n186# gnd 0.011519f
C68 a_270_n382# p3 0.060798f
C69 a_617_285# gnd 0.087075f
C70 a_594_556# p2 0.013746f
C71 a_617_285# a_600_239# 0.001275f
C72 w_417_462# a_397_472# 0.028268f
C73 w_259_n385# vdd 0.008451f
C74 g0 a_582_25# 0.003752f
C75 w_830_114# s1 0.013216f
C76 a_303_n248# gnd 0.396612f
C77 w_726_513# vdd 0.013119f
C78 g3 b3 0.756931f
C79 a_731_424# a_740_401# 0.001268f
C80 a_705_n209# p3 0.060798f
C81 p2 vdd 1.094079f
C82 w_611_305# a_617_318# 0.009864f
C83 a_825_350# gnd 0.247451f
C84 w_439_167# g0 4.29e-19
C85 w_538_625# vdd 0.008451f
C86 w_725_n171# p3 0.028748f
C87 w_401_n240# vdd 0.0086f
C88 w_238_456# a_251_466# 0.019526f
C89 g0 a0 0.001371f
C90 a_381_614# p2 0.005763f
C91 w_328_18# a_337_67# 0.027662f
C92 w_602_63# a_582_25# 0.026794f
C93 a_738_n161# vdd 0.019283f
C94 w_417_462# vdd 0.008451f
C95 w_676_271# c2 0.013216f
C96 a_380_291# p1g0 0.060798f
C97 a_743_378# gnd 0.247451f
C98 p1 a_269_n114# 0.060798f
C99 a_714_378# p2p1p0c0 7.68e-20
C100 w_226_594# vdd 6.13e-19
C101 a_610_395# p1 0.013746f
C102 w_764_n163# c3 1.23e-19
C103 w_720_n37# vdd 6.13e-19
C104 w_760_117# a_769_115# 0.027662f
C105 a_302_n114# gnd 0.396612f
C106 a_345_n42# vdd 0.439891f
C107 w_328_18# a_302_20# 0.007992f
C108 w_721_109# a_734_119# 0.015055f
C109 a_303_n248# a_338_n201# 0.063232f
C110 w_774_654# vdd 0.008451f
C111 a_397_472# a_440_412# 0.41238f
C112 w_302_599# a_239_604# 0.026907f
C113 w_400_323# a_380_291# 0.026907f
C114 a_440_393# gnd 0.41238f
C115 b0 a_582_25# 0.00288f
C116 w_877_383# p3p2p1p0c0 0.043313f
C117 a_883_389# p3p2p1g0 0.004158f
C118 a_302_20# a_345_92# 0.20619f
C119 w_807_654# cin 0.026794f
C120 w_258_n117# vdd 0.008451f
C121 a_733_n27# vdd 0.019283f
C122 w_726_513# g2 0.036563f
C123 a_731_492# a_731_457# 0.41238f
C124 a2 a_303_n248# 0.413834f
C125 a_518_635# g0 0.059018f
C126 a_883_429# p3p2p1g0 4.37e-21
C127 a_724_454# p2p1p0c0 2.55e-19
C128 a_445_147# a_490_101# 0.029681f
C129 a0 b0 0.704486f
C130 a_610_414# cin 0.013746f
C131 w_329_n250# b2 1.23e-19
C132 w_259_n251# a_270_n248# 0.026907f
C133 w_368_n246# a2 0.028748f
C134 w_400_28# vdd 0.0086f
C135 w_439_167# pocin 0.036563f
C136 a_457_101# gnd 0.247451f
C137 p1 a_769_115# 0.014473f
C138 g0 p2 0.010111f
C139 p3g2 gnd 0.207724f
C140 w_226_594# g2 0.008451f
C141 w_400_185# vdd 0.008451f
C142 c2 a_781_n52# 0.003948f
C143 a_734_119# gnd 0.396612f
C144 a_315_567# p3g2 0.060798f
C145 a_810_82# vdd 0.441416f
C146 a_251_466# gnd 0.701773f
C147 a_884_498# vdd 0.41238f
C148 w_725_444# a_724_454# 0.036563f
C149 a_883_396# a_825_350# 0.001275f
C150 w_725_266# vdd 0.0086f
C151 gnd p1g0 0.20619f
C152 w_687_n43# a_700_n75# 0.013216f
C153 w_758_272# cin 0.013592f
C154 a_594_575# a_594_556# 0.41238f
C155 a_819_257# gnd 0.011519f
C156 a_600_239# p1g0 7.68e-20
C157 w_797_280# p0 0.007896f
C158 a_380_153# vdd 0.441416f
C159 cin a_271_142# 0.001372f
C160 w_878_485# p3g2 0.036563f
C161 a_797_547# p3 0.013746f
C162 w_440_301# vdd 0.008451f
C163 w_796_n32# a_733_n27# 0.027261f
C164 w_599_n75# b1 0.009938f
C165 a_346_n310# vdd 0.439891f
C166 p2g1 a_776_378# 0.013746f
C167 w_367_n112# a_302_n114# 0.015055f
C168 p3 gnd 1.53153f
C169 w_472_604# p3p2g1 0.013216f
C170 a_738_234# gnd 0.20619f
C171 w_867_277# a_847_245# 0.026907f
C172 s0 vdd 0.439883f
C173 a1 a_302_n114# 0.413834f
C174 w_620_464# a_534_474# 0.028268f
C175 p0 cin 0.001461f
C176 a_688_664# vdd 2.20188f
C177 s3 gnd 0.20619f
C178 a_270_n382# a_303_n382# 0.060798f
C179 a_440_412# g0 0.013746f
C180 b3 a_346_n310# 0.012282f
C181 a3 a_582_n389# 0.060856f
C182 a_731_424# a_743_378# 0.002189f
C183 w_725_411# p2p1p0c0 0.001078f
C184 a_617_285# vdd 0.001532f
C185 a_847_245# gnd 0.248155f
C186 w_384_462# a_397_472# 0.018373f
C187 g0 a_490_101# 0.013746f
C188 w_834_n166# vdd 0.008451f
C189 a_453_311# p1 0.002443f
C190 a_424_554# p2 0.013746f
C191 a_303_n248# vdd 0.019283f
C192 w_658_464# vdd 0.008451f
C193 a_270_n248# gnd 0.248155f
C194 g3 a3 0.001371f
C195 a_883_429# a_883_389# 0.41238f
C196 w_611_340# a_617_318# 0.009864f
C197 a_892_373# p3p2p1g0 2.36e-20
C198 w_505_625# vdd 0.008451f
C199 a_617_285# p1p0c0 0.192837f
C200 w_368_n246# vdd 6.13e-19
C201 w_692_n177# p3 0.028034f
C202 w_569_57# a_582_25# 0.013216f
C203 a_773_n165# vdd 9.08e-21
C204 a_781_n52# gnd 0.011519f
C205 w_384_462# vdd 0.008451f
C206 w_879_518# g3 0.036563f
C207 a_705_n209# c3 1.47e-20
C208 a_731_424# a_731_417# 0.453641f
C209 p3g2 a_883_396# 0.001345f
C210 a_714_378# gnd 0.247451f
C211 a_302_20# a_337_67# 0.063232f
C212 w_193_588# vdd 0.0086f
C213 w_368_604# p3 0.026794f
C214 w_725_n171# c3 0.013592f
C215 w_687_n43# vdd 0.0086f
C216 a_806_278# a_771_282# 0.063232f
C217 w_400_28# b0 0.015139f
C218 w_569_57# a0 0.028093f
C219 w_291_17# a_302_20# 0.027261f
C220 a_302_n114# vdd 0.019283f
C221 w_741_654# vdd 0.008451f
C222 w_642_625# p3p2p1g0 0.013216f
C223 a_594_575# g0 0.013746f
C224 w_760_117# p1 0.007896f
C225 a_269_n114# gnd 0.248155f
C226 w_226_594# a_239_604# 0.019526f
C227 a_734_119# c1 0.599413f
C228 w_367_323# a_380_291# 0.013216f
C229 a0 a_582_25# 0.060867f
C230 a_876_426# p3p2p1g0 2.55e-19
C231 w_401_n240# a_346_n176# 0.013216f
C232 w_830_114# vdd 0.008451f
C233 w_329_n250# a_338_n201# 0.027662f
C234 w_845_654# a_688_664# 0.027163f
C235 a_768_n31# vdd 9.08e-21
C236 a_782_94# gnd 0.011519f
C237 a_731_492# p2g1g0 3.63e-19
C238 b2 a_325_n180# 0.003948f
C239 p3p2g1 p3p2p1g0 0.00851f
C240 a_445_147# a_457_101# 0.001275f
C241 w_367_22# vdd 6.13e-19
C242 a_610_414# p0 0.013746f
C243 w_759_n29# p2 0.007896f
C244 w_329_n250# a2 0.007896f
C245 a_738_n161# a_814_n198# 0.060798f
C246 a_345_92# gnd 0.20619f
C247 w_400_185# pocin 0.013216f
C248 a_617_285# g1 1.39e-20
C249 p2p1g0 gnd 0.20619f
C250 p3g2 vdd 0.440124f
C251 w_367_185# vdd 0.008507f
C252 a_734_119# vdd 0.019283f
C253 w_790_410# a_731_424# 0.027289f
C254 a_380_153# pocin 0.060798f
C255 a_424_535# gnd 0.41238f
C256 a_251_466# vdd 0.017997f
C257 w_676_271# vdd 0.008451f
C258 vdd p1g0 0.439883f
C259 gnd p3p2p1g0 0.20619f
C260 a_662_239# gnd 0.247451f
C261 w_758_272# p0 0.028748f
C262 a_302_n114# a_337_n67# 0.063232f
C263 p0 a_271_142# 0.060798f
C264 w_328_n116# a_302_n114# 0.007992f
C265 w_400_323# vdd 0.008451f
C266 a_610_395# a_610_377# 0.41238f
C267 a_303_n382# gnd 0.396612f
C268 w_759_n29# a_733_n27# 0.007992f
C269 p3 vdd 1.414045f
C270 w_834_277# a_847_245# 0.013216f
C271 w_473_301# p0 0.026996f
C272 a_304_190# gnd 0.701773f
C273 a_738_234# vdd 0.439891f
C274 b1 a_324_n46# 0.003948f
C275 w_726_513# a_731_492# 0.009864f
C276 a_381_614# p3 0.002443f
C277 w_587_464# a_534_474# 0.028268f
C278 w_879_518# a_884_498# 0.009864f
C279 a3 a_346_n310# 0.060798f
C280 g3 a_582_n389# 0.003752f
C281 s3 vdd 0.439883f
C282 w_790_410# vdd 0.008451f
C283 w_725_444# p2p1p0c0 2.18e-19
C284 a_688_664# cin 0.059018f
C285 a_325_n314# a_303_n382# 0.080021f
C286 c3 gnd 0.20621f
C287 a_731_424# a_714_378# 0.002189f
C288 w_335_599# p3g2 0.013216f
C289 w_554_464# p1 0.026794f
C290 a_733_n27# a_809_n64# 0.060798f
C291 a_847_245# vdd 0.441416f
C292 a_771_282# gnd 0.396612f
C293 w_602_n351# b3 0.008451f
C294 w_801_n166# vdd 0.008507f
C295 w_238_456# a_218_418# 0.026794f
C296 w_368_n380# a_303_n382# 0.015055f
C297 a_797_566# p2 0.013746f
C298 a_325_n180# gnd 0.011519f
C299 w_620_464# vdd 0.008451f
C300 a_270_n248# vdd 0.441416f
C301 a_731_417# p2g1 0.015843f
C302 a_617_318# vdd 0.41238f
C303 a_453_311# gnd 0.042086f
C304 c1 a_782_94# 0.003948f
C305 w_472_604# vdd 0.008451f
C306 w_329_n250# vdd 0.001288f
C307 a_617_285# a_617_278# 0.453641f
C308 a_518_635# p2 0.004034f
C309 w_347_461# vdd 0.008451f
C310 s2 gnd 0.20619f
C311 a_731_457# a_731_417# 0.41238f
C312 w_538_625# a_518_635# 0.028268f
C313 w_472_604# a_381_614# 0.027163f
C314 a_693_378# gnd 0.247451f
C315 g0 p1g0 0.007385f
C316 a_251_466# g1 0.740337f
C317 a_453_311# a_496_251# 0.41238f
C318 a_324_n46# gnd 0.011519f
C319 g1 p1g0 0.00851f
C320 w_708_654# vdd 0.008451f
C321 a_688_664# p3p2p1p0c0 0.060798f
C322 w_721_109# p1 0.028748f
C323 w_400_28# a0 0.028034f
C324 w_291_17# a_269_20# 0.013216f
C325 w_367_22# b0 0.014021f
C326 a_303_n248# a_346_n176# 0.20619f
C327 a_269_n114# vdd 0.441416f
C328 w_400_323# g0 0.011382f
C329 a_883_396# p3p2p1g0 0.040586f
C330 a_269_20# a_302_20# 0.060798f
C331 w_774_654# p0 0.026996f
C332 a_769_115# c1 5.8e-19
C333 a_734_119# a_701_71# 0.20619f
C334 w_538_625# p2 0.026794f
C335 w_807_654# a_688_664# 0.028268f
C336 w_834_n166# a_814_n198# 0.026907f
C337 w_797_114# vdd 0.008507f
C338 a_397_472# p2p1g0 0.060798f
C339 w_720_n37# p2 0.028748f
C340 w_328_18# vdd 0.001288f
C341 a_534_474# p1 0.004034f
C342 a_251_466# a_327_429# 0.060798f
C343 a_302_20# gnd 0.396612f
C344 a_345_92# vdd 0.439891f
C345 a_218_418# gnd 0.20619f
C346 a_534_474# p2p1p0c0 0.060798f
C347 p2p1g0 vdd 0.439883f
C348 w_829_n32# s2 0.013216f
C349 w_291_180# vdd 6.13e-19
C350 p1 gnd 0.684683f
C351 a_769_115# vdd 9.08e-21
C352 a_733_n27# p2 0.413834f
C353 w_725_411# a_731_424# 0.013329f
C354 a_594_537# gnd 0.41238f
C355 a_731_424# c3 0.060798f
C356 vdd p3p2p1g0 0.439883f
C357 gnd p2p1p0c0 0.20619f
C358 w_258_312# p1 0.028034f
C359 w_725_266# p0 0.028034f
C360 a_629_239# gnd 0.247451f
C361 w_347_461# p2g1 0.013216f
C362 a_206_556# gnd 0.20619f
C363 cin a_819_257# 0.003948f
C364 w_759_n29# a_768_n31# 0.027662f
C365 w_599_n75# g1 0.019526f
C366 w_720_n37# a_733_n27# 0.015055f
C367 w_400_n106# b1 0.015139f
C368 w_566_n81# a1 0.028089f
C369 w_291_n117# a_302_n114# 0.027261f
C370 w_367_323# vdd 0.008493f
C371 a_303_n382# vdd 0.019283f
C372 a_270_n382# gnd 0.248155f
C373 a_518_635# a_594_575# 0.41238f
C374 w_834_277# a_771_282# 0.027261f
C375 a_626_262# gnd 0.001534f
C376 w_611_272# p1p0c0 0.043313f
C377 a_617_278# p1g0 0.004158f
C378 a_304_190# vdd 0.017997f
C379 w_488_462# p2p1g0 0.013216f
C380 a_239_604# p3 0.001371f
C381 p1p0c0 a_662_239# 0.013746f
C382 a_738_234# cin 1.47e-20
C383 w_569_n357# vdd 0.008451f
C384 w_554_464# a_534_474# 0.028268f
C385 a_705_n209# gnd 0.20619f
C386 b3 a_303_n382# 0.599413f
C387 c3 vdd 0.439883f
C388 a_731_424# a_693_378# 0.001275f
C389 a_883_396# a_883_389# 0.453641f
C390 a_688_664# p0 0.005763f
C391 a_771_282# vdd 0.019283f
C392 a_271_280# p1 0.060798f
C393 w_347_461# a_327_429# 0.026907f
C394 w_764_n163# vdd 0.001288f
C395 w_205_450# a_218_418# 0.013216f
C396 w_329_n384# a_303_n382# 0.007992f
C397 w_760_117# c1 1.23e-19
C398 b2 gnd 0.037678f
C399 w_587_464# vdd 0.008451f
C400 a_892_373# gnd 0.001534f
C401 w_544_301# a_453_311# 0.027163f
C402 w_620_464# cin 0.026794f
C403 a_453_311# vdd 1.32165f
C404 w_434_604# vdd 0.008451f
C405 a_610_377# p1 0.013746f
C406 w_292_n251# vdd 0.008507f
C407 a_688_664# p2 0.004034f
C408 w_314_461# vdd 0.008507f
C409 c2 gnd 0.20621f
C410 s2 vdd 0.439883f
C411 w_434_604# a_381_614# 0.028268f
C412 w_505_625# a_518_635# 0.018373f
C413 a_380_291# gnd 0.248155f
C414 w_291_318# a_271_280# 0.026794f
C415 w_566_n81# vdd 0.008451f
C416 a_453_311# p1p0c0 0.060798f
C417 a_617_318# a_617_278# 0.41238f
C418 w_692_n177# a_705_n209# 0.013216f
C419 w_571_625# p1 0.026996f
C420 w_328_18# b0 1.23e-19
C421 w_688_103# p1 0.028034f
C422 w_258_17# a_269_20# 0.026907f
C423 w_367_22# a0 0.028748f
C424 b2 a_338_n201# 5.8e-19
C425 w_675_654# vdd 0.008451f
C426 b1 gnd 0.036517f
C427 a_738_n161# a_786_n186# 0.080021f
C428 a_814_n198# s3 0.060798f
C429 b0 a_345_92# 0.012282f
C430 a_324_88# a_302_20# 0.080021f
C431 p1 c1 0.001461f
C432 w_367_323# g0 0.011382f
C433 w_760_117# vdd 0.001288f
C434 w_801_n166# a_814_n198# 0.013216f
C435 w_774_654# a_688_664# 0.028268f
C436 a2 b2 0.696062f
C437 w_384_462# p2 0.026794f
C438 a_884_498# a_883_464# 0.41238f
C439 a_337_67# vdd 9.08e-21
C440 s1 gnd 0.20619f
C441 a_731_424# p2p1p0c0 0.040586f
C442 p3p2g1 gnd 0.207724f
C443 w_291_17# vdd 0.008507f
C444 w_687_n43# p2 0.028034f
C445 a_397_472# p1 0.005763f
C446 w_604_625# vdd 0.008451f
C447 a_269_20# gnd 0.248155f
C448 a_302_20# vdd 0.019283f
C449 w_400_185# a_380_153# 0.026907f
C450 a_773_n165# a_738_n161# 0.063232f
C451 a_218_418# vdd 0.439891f
C452 a_534_474# gnd 0.042086f
C453 a_440_393# p2 0.013746f
C454 w_725_411# p2g1 0.043313f
C455 w_258_174# vdd 0.0086f
C456 a_594_556# p1 0.013746f
C457 a_424_554# a_424_535# 0.41238f
C458 a_768_n31# p2 0.014473f
C459 a_700_n75# c2 1.47e-20
C460 a_594_556# a_594_537# 0.41238f
C461 w_291_180# cin 0.008451f
C462 p1 vdd 0.681699f
C463 w_877_451# a_883_464# 0.01128f
C464 a_797_547# gnd 0.41238f
C465 a_496_232# p1 0.013746f
C466 w_434_604# g1 0.026794f
C467 a_883_396# a_892_373# 0.001268f
C468 w_611_340# gnd 9.65e-20
C469 vdd p2p1p0c0 0.439883f
C470 w_599_n75# a_579_n113# 0.026794f
C471 a_797_585# a_797_566# 0.41238f
C472 a_302_n114# a_345_n42# 0.20619f
C473 a_600_239# gnd 0.247451f
C474 a_315_567# gnd 0.248155f
C475 a_206_556# vdd 0.439891f
C476 a_797_604# cin 0.013746f
C477 w_400_n106# a1 0.028034f
C478 w_291_n117# a_269_n114# 0.013216f
C479 w_367_n112# b1 0.014021f
C480 a_303_n382# a_338_n335# 0.063232f
C481 a_270_n382# vdd 0.441416f
C482 w_877_383# p3p2p1g0 0.001078f
C483 a_797_585# p0 0.013746f
C484 w_291_318# vdd 6.13e-19
C485 a_325_n314# gnd 0.011519f
C486 a_610_315# p1g0 2.55e-19
C487 a1 b1 0.779908f
C488 w_611_272# a_617_278# 0.017071f
C489 w_797_280# a_771_282# 0.007992f
C490 w_401_n374# vdd 0.0086f
C491 a_518_635# p3 0.002443f
C492 a_251_466# p2 0.001371f
C493 a_738_234# p0 0.060798f
C494 w_602_n351# a_582_n389# 0.026794f
C495 w_521_464# a_534_474# 0.018373f
C496 a_304_190# cin 0.740337f
C497 a_610_414# a_610_395# 0.41238f
C498 a_705_n209# vdd 0.439891f
C499 a3 a_303_n382# 0.413834f
C500 a_440_412# a_440_393# 0.41238f
C501 a_866_350# p3p2p1g0 7.68e-20
C502 a_768_n31# a_733_n27# 0.063232f
C503 a_928_350# gnd 0.247451f
C504 a_806_278# vdd 9.08e-21
C505 w_604_625# g0 0.026794f
C506 a_771_282# cin 0.599413f
C507 w_401_n374# b3 0.015139f
C508 w_292_n385# a_303_n382# 0.027261f
C509 w_259_n385# p3 0.013216f
C510 w_314_461# a_327_429# 0.013216f
C511 w_569_n357# a3 0.02808f
C512 w_602_n351# g3 0.019526f
C513 w_725_n171# vdd 6.13e-19
C514 w_554_464# vdd 0.008451f
C515 g2 p2p1p0c0 0.054984f
C516 p3p2g1 a_883_396# 0.001345f
C517 w_721_109# c1 0.013592f
C518 b2 vdd 2.33e-19
C519 a2 gnd 1.559369f
C520 w_726_513# p3 4.5e-19
C521 a_271_280# gnd 0.20619f
C522 w_506_301# a_453_311# 0.028268f
C523 w_401_604# vdd 0.008451f
C524 w_259_n251# vdd 0.008451f
C525 a_218_418# g1 0.001372f
C526 a_206_556# g2 0.001372f
C527 g0 p1 0.015049f
C528 a_453_311# cin 0.059018f
C529 a_738_n161# p3 0.413834f
C530 w_830_114# a_810_82# 0.026907f
C531 a_700_n75# gnd 0.20619f
C532 c2 vdd 0.439883f
C533 w_238_456# vdd 6.13e-19
C534 w_401_604# a_381_614# 0.028268f
C535 b0 a_337_67# 5.8e-19
C536 a_380_291# vdd 0.441416f
C537 w_258_312# a_271_280# 0.013216f
C538 a_610_377# gnd 0.41238f
C539 w_400_n106# vdd 0.0086f
C540 a_270_n248# p2 0.060798f
C541 w_328_18# a0 0.007896f
C542 a1 gnd 1.537765f
C543 b2 a_582_n251# 0.002958f
C544 a2 a_338_n201# 0.014473f
C545 b1 vdd 2.33e-19
C546 w_642_625# vdd 0.008451f
C547 w_291_318# g0 0.008451f
C548 w_367_323# a_304_328# 0.026907f
C549 a_883_396# gnd 0.099139f
C550 b0 a_302_20# 0.599413f
C551 a0 a_345_92# 0.060798f
C552 p1 a_701_71# 0.060798f
C553 w_721_109# vdd 6.13e-19
C554 w_741_654# a_688_664# 0.028268f
C555 w_368_n246# a_303_n248# 0.015055f
C556 a_610_395# p0 0.013746f
C557 w_801_n166# a_738_n161# 0.027261f
C558 w_602_n213# b2 0.008451f
C559 a_884_498# p3g2 3.63e-19
C560 c1 gnd 0.20621f
C561 s1 vdd 0.439883f
C562 g2 b2 0.757544f
C563 a_734_119# a_810_82# 0.060798f
C564 w_877_383# a_883_389# 0.017071f
C565 p3p2g1 vdd 0.439963f
C566 a_731_424# gnd 0.093107f
C567 a_731_457# p2p1p0c0 4.37e-21
C568 w_258_17# vdd 0.008451f
C569 w_708_654# p2 0.026794f
C570 w_291_180# a_271_142# 0.026794f
C571 w_367_185# a_380_153# 0.013216f
C572 a_324_88# gnd 0.011519f
C573 a_269_20# vdd 0.441416f
C574 a_381_614# p3p2g1 0.060798f
C575 a_397_472# gnd 0.042086f
C576 a_534_474# vdd 1.76176f
C577 a_445_147# a_445_140# 0.453641f
C578 w_867_277# vdd 0.008451f
C579 a_883_396# a_928_350# 0.029681f
C580 a_445_140# vdd 0.41238f
C581 a_445_147# gnd 0.081043f
C582 w_725_444# a_731_457# 0.009864f
C583 g0 a_380_291# 0.008577f
C584 a_883_389# p3p2p1p0c0 0.015843f
C585 w_566_n81# a_579_n113# 0.013216f
C586 vdd gnd 2.215758f
C587 w_611_340# vdd 0.013119f
C588 w_725_266# a_738_234# 0.013216f
C589 w_238_456# g1 0.008451f
C590 b1 a_337_n67# 5.8e-19
C591 a_496_232# gnd 0.41238f
C592 a_733_n27# a_781_n52# 0.080021f
C593 a_809_n64# s2 0.060798f
C594 a_518_635# p3p2p1g0 0.060798f
C595 a_381_614# gnd 0.042086f
C596 a_304_190# a_271_142# 0.003752f
C597 a_315_567# vdd 0.441416f
C598 w_877_416# p3p2p1g0 2.18e-19
C599 w_258_312# vdd 0.0086f
C600 b3 gnd 0.03396f
C601 a_797_604# p0 0.013746f
C602 w_328_n116# b1 1.23e-19
C603 w_258_n117# a_269_n114# 0.026907f
C604 w_367_n112# a1 0.028748f
C605 g1 b1 0.7623f
C606 w_797_280# a_806_278# 0.027662f
C607 w_676_271# a_617_285# 0.027289f
C608 w_611_305# a_617_278# 0.008113f
C609 w_758_272# a_771_282# 0.015055f
C610 a_239_604# a_206_556# 0.003752f
C611 a_617_285# p1g0 0.040586f
C612 p1p0c0 gnd 0.207724f
C613 w_569_n357# a_582_n389# 0.013216f
C614 a_688_664# p3 0.002443f
C615 a_424_535# p2 0.013746f
C616 a_496_251# a_496_232# 0.41238f
C617 a_304_190# p0 0.001371f
C618 w_368_n380# vdd 6.13e-19
C619 a_338_n201# vdd 9.08e-21
C620 b3 a_325_n314# 0.003948f
C621 a_582_n251# gnd 0.20619f
C622 a_895_350# gnd 0.247451f
C623 a_847_245# s0 0.060798f
C624 a_771_282# p0 0.413834f
C625 w_692_n177# vdd 0.0086f
C626 a_806_278# cin 5.8e-19
C627 w_401_n374# a3 0.028034f
C628 w_292_n385# a_270_n382# 0.013216f
C629 w_368_n380# b3 0.014021f
C630 a2 vdd 0.228122f
C631 c3 g3 0.054984f
C632 g2 gnd 0.661342f
C633 w_521_464# vdd 0.008451f
C634 c4 gnd 0.20619f
C635 a_271_280# vdd 0.439891f
C636 w_473_301# a_453_311# 0.028268f
C637 w_587_464# p0 0.026996f
C638 w_368_604# vdd 0.008451f
C639 w_505_625# p3 0.026794f
C640 g0 a_445_140# 0.016231f
C641 w_834_n166# s3 0.013216f
C642 a_453_311# p0 0.005763f
C643 a_304_328# p1 0.001371f
C644 w_829_n32# vdd 0.008451f
C645 w_205_450# vdd 0.0086f
C646 w_400_28# a_345_92# 0.013216f
C647 w_504_133# c1 0.013216f
C648 a_773_n165# p3 0.014473f
C649 a_700_n75# vdd 0.439891f
C650 w_797_114# a_810_82# 0.013216f
C651 w_368_604# a_381_614# 0.018373f
C652 w_335_599# a_315_567# 0.026907f
C653 g0 gnd 0.207724f
C654 a0 a_337_67# 0.014473f
C655 w_193_588# p3 0.028034f
C656 w_367_n112# vdd 6.13e-19
C657 b2 a_346_n176# 0.012282f
C658 a2 a_582_n251# 0.060856f
C659 a_270_n248# a_303_n248# 0.060798f
C660 w_611_340# g1 0.036563f
C661 a1 vdd 0.228122f
C662 a_738_n161# c3 0.599413f
C663 g1 gnd 0.661342f
C664 a0 a_302_20# 0.413834f
C665 p2g1 gnd 0.207724f
C666 a_883_396# vdd 0.001532f
C667 w_291_318# a_304_328# 0.019526f
C668 a_445_147# c1 0.060798f
C669 w_571_625# vdd 0.008451f
C670 w_329_n250# a_303_n248# 0.007992f
C671 w_708_654# a_688_664# 0.028268f
C672 w_764_n163# a_738_n161# 0.007992f
C673 w_688_103# vdd 0.0086f
C674 g2 a2 0.001371f
C675 c1 vdd 0.439883f
C676 w_504_133# a_445_147# 0.027289f
C677 w_439_134# a_445_140# 0.017071f
C678 a_701_71# gnd 0.20619f
C679 a_731_424# vdd 0.001532f
C680 p2g1g0 p2p1p0c0 0.00851f
C681 w_942_382# a_883_396# 0.027289f
C682 w_877_416# a_883_389# 0.008113f
C683 w_504_133# vdd 0.008451f
C684 w_258_174# a_271_142# 0.013216f
C685 b0 gnd 0.035313f
C686 pocin a_445_140# 0.185571f
C687 w_877_416# a_883_429# 0.009864f
C688 a_327_429# gnd 0.248155f
C689 a_397_472# vdd 1.32165f
C690 w_604_625# a_518_635# 0.028268f
C691 w_834_277# vdd 0.008507f
C692 a_797_566# p1 0.013746f
C693 w_759_n29# c2 1.23e-19
C694 a_883_396# a_895_350# 0.002189f
C695 g0 a_271_280# 0.001372f
C696 a_534_474# cin 0.059018f
C697 pocin gnd 0.372676f
C698 a_445_147# vdd 0.001532f
C699 w_258_174# p0 0.028034f
C700 w_544_301# vdd 0.008451f
C701 w_400_323# p1g0 0.013216f
C702 a_518_635# p1 0.005763f
C703 a_883_396# c4 0.060798f
C704 a_304_328# a_380_291# 0.060798f
C705 a_269_n114# a_302_n114# 0.060798f
C706 cin gnd 1.99e-20
C707 b1 a_579_n113# 0.00343f
C708 a1 a_337_n67# 0.014473f
C709 a_381_614# vdd 1.32165f
C710 a_239_604# gnd 0.248155f
C711 a_304_190# a_380_153# 0.060798f
C712 a_218_418# p2 0.060798f
C713 a_731_424# g2 1.39e-20
C714 w_328_n116# a1 0.007896f
C715 b3 vdd 2.33e-19
C716 a_303_n382# a_346_n310# 0.20619f
C717 w_942_382# vdd 0.008451f
C718 a3 gnd 0.414526f
C719 p1p0c0 vdd 0.439883f
C720 w_544_301# p1p0c0 0.013216f
C721 a_688_664# a_797_604# 0.41238f
C722 g1 a1 0.001371f
C723 w_611_305# a_610_315# 0.036563f
C724 w_611_272# a_617_285# 0.013329f
C725 a_239_604# a_315_567# 0.060798f
C726 w_329_n384# vdd 0.001288f
C727 a_594_537# p2 0.013746f
C728 g0 c1 0.008006f
C729 w_488_462# a_397_472# 0.027163f
C730 a_617_285# a_662_239# 0.029681f
C731 a_496_251# cin 0.013746f
C732 a_582_n251# vdd 0.439883f
C733 a_346_n176# gnd 0.20619f
C734 w_504_133# g0 0.011197f
C735 a_866_350# gnd 0.247451f
C736 w_417_462# p1 0.026996f
C737 a_617_318# p1g0 4.37e-21
C738 w_329_n384# b3 1.23e-19
C739 w_259_n385# a_270_n382# 0.026907f
C740 w_368_n380# a3 0.028748f
C741 a_806_278# p0 0.014473f
C742 c3 a_786_n186# 0.003948f
C743 w_688_103# a_701_71# 0.013216f
C744 w_488_462# vdd 0.008451f
C745 a_397_472# g0 0.059018f
C746 a_731_424# p2g1 0.192837f
C747 a_814_n198# gnd 0.248155f
C748 g2 vdd 0.022667f
C749 a_701_71# c1 1.47e-20
C750 p3p2p1p0c0 gnd 0.207724f
C751 w_440_301# a_453_311# 0.018373f
C752 c4 vdd 0.439883f
C753 w_335_599# vdd 0.008451f
C754 g0 a_445_147# 0.202944f
C755 w_796_n32# vdd 0.008507f
C756 w_797_114# a_734_119# 0.027261f
C757 a_579_n113# gnd 0.20619f
C758 a_337_n67# vdd 9.08e-21
C759 a_883_464# a_883_429# 0.41238f
C760 a_534_474# a_610_414# 0.41238f
C761 w_258_n117# p1 0.013216f
C762 w_845_654# vdd 0.008451f
C763 w_226_594# a_206_556# 0.026794f
C764 w_302_599# a_315_567# 0.013216f
C765 a_734_119# a_782_94# 0.080021f
C766 w_544_301# g0 0.00229f
C767 w_942_382# c4 0.013216f
C768 a_740_401# p2p1p0c0 2.36e-20
C769 g0 vdd 0.122827f
C770 a_304_328# gnd 0.701773f
C771 w_328_n116# vdd 0.001288f
C772 w_602_n213# a_582_n251# 0.026794f
C773 a_440_412# p1 0.013746f
C774 a_325_n180# a_303_n248# 0.080021f
C775 a_773_n165# c3 5.8e-19
C776 a_738_n161# a_705_n209# 0.20619f
C777 a2 a_346_n176# 0.060798f
C778 g2 a_582_n251# 0.003752f
C779 a_809_n64# gnd 0.248155f
C780 g1 vdd 0.024039f
C781 p2g1 vdd 0.439883f
C782 b0 a_324_88# 0.003948f
C783 w_401_604# p2 0.026996f
C784 g0 p1p0c0 0.002352f
C785 p3p2p1p0c0 a_928_350# 0.013746f
C786 a_381_614# g1 0.059018f
C787 w_292_n251# a_303_n248# 0.027261f
C788 w_259_n251# p2 0.013216f
C789 w_675_654# a_688_664# 0.018373f
C790 w_642_625# a_518_635# 0.027163f
C791 w_401_n240# b2 0.015139f
C792 w_764_n163# a_773_n165# 0.027662f
C793 w_569_n219# a2 0.028079f
C794 w_602_n213# g2 0.019526f
C795 w_725_n171# a_738_n161# 0.015055f
C796 w_439_167# a_445_140# 0.008113f
C797 w_439_134# a_445_147# 0.013329f
C798 a_582_25# gnd 0.20619f
C799 a_701_71# vdd 0.439891f
C800 c2 p2 0.001461f
C801 a_769_115# a_734_119# 0.063232f
C802 w_877_416# a_876_426# 0.036563f
C803 w_877_383# a_883_396# 0.013329f
C804 p2g1g0 gnd 0.001534f
C805 w_258_17# p0 0.013216f
C806 a0 gnd 1.211792f
C807 b0 vdd 2.33e-19
C808 w_725_411# a_731_417# 0.017071f
C809 pocin a_445_147# 1.39e-20
C810 p0 a_269_20# 0.060798f
C811 a_327_429# vdd 0.441416f
C812 w_877_451# a_883_429# 0.009864f
C813 a_883_396# a_866_350# 0.002189f
C814 a_534_474# p0 0.005763f
C815 w_797_280# vdd 0.001288f
C816 a_304_328# a_271_280# 0.003752f
C817 w_611_272# p1g0 0.001078f
C818 a_594_575# p1 0.013746f
C819 w_720_n37# c2 0.013592f
C820 w_440_301# p1 0.026794f
C821 w_367_185# a_304_190# 0.026907f
C822 a_797_566# a_797_547# 0.41238f
C823 pocin vdd 0.439883f
C824 a_271_142# gnd 0.20619f
C825 w_725_479# a_731_457# 0.009864f
C826 a_424_535# p3 0.013746f
C827 a_582_n389# gnd 0.20619f
C828 a_883_396# p3p2p1p0c0 0.192837f
C829 a_688_664# p1 0.004034f
C830 w_506_301# vdd 0.008451f
C831 w_829_n32# a_809_n64# 0.026907f
C832 w_328_n116# a_337_n67# 0.027662f
C833 w_400_n106# a_345_n42# 0.013216f
C834 a_338_n335# vdd 9.08e-21
C835 b1 a_345_n42# 0.012282f
C836 a1 a_579_n113# 0.060856f
C837 a_797_604# a_797_585# 0.41238f
C838 cin vdd 0.024438f
C839 a_324_n46# a_302_n114# 0.080021f
C840 a_733_n27# c2 0.599413f
C841 a_381_614# a_424_554# 0.41238f
C842 p0 gnd 0.628007f
C843 a_534_474# p2 0.002443f
C844 a_518_635# gnd 0.042086f
C845 a_239_604# vdd 0.017997f
C846 g3 gnd 0.661342f
C847 b3 a_338_n335# 5.8e-19
C848 a3 vdd 0.228122f
C849 w_602_63# g0 0.019526f
C850 w_450_462# a_397_472# 0.028268f
C851 a_617_285# a_629_239# 0.002189f
C852 a_771_282# a_819_257# 0.080021f
C853 a_797_547# p2 0.013746f
C854 a_496_251# p0 0.013746f
C855 w_329_n384# a_338_n335# 0.027662f
C856 w_401_n374# a_346_n310# 0.013216f
C857 w_292_n385# vdd 0.008507f
C858 w_879_518# vdd 0.013167f
C859 c3 p3 0.001461f
C860 p2 gnd 0.699156f
C861 a_346_n176# vdd 0.439891f
C862 w_658_464# p2p1p0c0 0.013216f
C863 a3 b3 0.700527f
C864 w_439_134# g0 0.051169f
C865 a_845_350# gnd 0.247451f
C866 w_764_n163# p3 0.007896f
C867 a_617_285# a_626_262# 0.001268f
C868 a_617_278# p1p0c0 0.015843f
C869 w_314_461# a_251_466# 0.026907f
C870 g0 b0 0.756776f
C871 w_329_n384# a3 0.007896f
C872 a_771_282# a_738_234# 0.20619f
C873 w_569_n219# vdd 0.008451f
C874 a_814_n198# vdd 0.441416f
C875 w_790_410# c3 0.013216f
C876 a_738_n161# gnd 0.396612f
C877 w_450_462# vdd 0.008451f
C878 p3p2p1p0c0 vdd 0.439883f
C879 w_741_654# p1 0.026794f
C880 a_776_378# gnd 0.247451f
C881 w_302_599# vdd 0.008507f
C882 a_771_282# a_847_245# 0.060798f
C883 w_759_n29# vdd 0.001288f
C884 a_239_604# g2 0.740337f
C885 a_440_393# p1 0.013746f
C886 w_367_22# a_302_20# 0.015055f
C887 w_602_63# b0 0.008938f
C888 a_883_464# p3p2g1 3.63e-19
C889 p2g1g0 a_731_424# 0.001345f
C890 a_327_429# p2g1 0.060798f
C891 a_345_n42# gnd 0.20619f
C892 w_807_654# vdd 0.008451f
C893 a_579_n113# vdd 0.439883f
C894 w_760_117# a_734_119# 0.007992f
C895 w_193_588# a_206_556# 0.013216f
C896 a_304_328# vdd 0.017767f
C897 a_810_82# s1 0.060798f
C898 a_740_401# gnd 0.001534f
C899 w_569_n219# a_582_n251# 0.013216f
C900 a_424_554# g1 0.013746f
C901 w_291_n117# vdd 0.008507f
C902 p1g0 0 1.041374f **FLOATING
C903 p3p2p1g0 0 1.051177f **FLOATING
C904 p2p1p0c0 0 1.047217f **FLOATING
C905 gnd 0 16.630608f **FLOATING
C906 vdd 0 29.946383f **FLOATING
C907 a_338_n335# 0 0.100202f **FLOATING
C908 a_582_n389# 0 0.477455f **FLOATING
C909 a_346_n310# 0 0.326258f **FLOATING
C910 p3 0 4.246335f **FLOATING
C911 a_303_n382# 0 0.665072f **FLOATING
C912 a_270_n382# 0 0.382299f **FLOATING
C913 a_325_n314# 0 0.12884f **FLOATING
C914 b3 0 6.48067f **FLOATING
C915 a3 0 2.52216f **FLOATING
C916 g3 0 1.415272f **FLOATING
C917 a_786_n186# 0 0.12884f **FLOATING
C918 s3 0 0.145867f **FLOATING
C919 c3 0 1.29723f **FLOATING
C920 a_705_n209# 0 0.326258f **FLOATING
C921 a_338_n201# 0 0.100202f **FLOATING
C922 a_582_n251# 0 0.477455f **FLOATING
C923 a_346_n176# 0 0.326258f **FLOATING
C924 p2 0 5.260555f **FLOATING
C925 a_303_n248# 0 0.665072f **FLOATING
C926 a_270_n248# 0 0.382299f **FLOATING
C927 a_325_n180# 0 0.12884f **FLOATING
C928 b2 0 6.40557f **FLOATING
C929 a2 0 2.41341f **FLOATING
C930 g2 0 1.459106f **FLOATING
C931 a_814_n198# 0 0.382299f **FLOATING
C932 a_738_n161# 0 0.665072f **FLOATING
C933 a_773_n165# 0 0.100202f **FLOATING
C934 a_781_n52# 0 0.12884f **FLOATING
C935 s2 0 0.145867f **FLOATING
C936 c2 0 1.30119f **FLOATING
C937 a_700_n75# 0 0.326258f **FLOATING
C938 a_337_n67# 0 0.100202f **FLOATING
C939 a_579_n113# 0 0.477455f **FLOATING
C940 a_345_n42# 0 0.326258f **FLOATING
C941 a_302_n114# 0 0.665072f **FLOATING
C942 a_269_n114# 0 0.382299f **FLOATING
C943 a_324_n46# 0 0.12884f **FLOATING
C944 b1 0 6.36751f **FLOATING
C945 a1 0 2.43873f **FLOATING
C946 g1 0 1.706117f **FLOATING
C947 a_809_n64# 0 0.382299f **FLOATING
C948 a_733_n27# 0 0.665072f **FLOATING
C949 a_768_n31# 0 0.100202f **FLOATING
C950 a_782_94# 0 0.12884f **FLOATING
C951 a_337_67# 0 0.100202f **FLOATING
C952 s1 0 0.145867f **FLOATING
C953 c1 0 1.30119f **FLOATING
C954 a_701_71# 0 0.326258f **FLOATING
C955 a_582_25# 0 0.477455f **FLOATING
C956 a_490_101# 0 0.019534f **FLOATING
C957 a_457_101# 0 0.024435f **FLOATING
C958 a_345_92# 0 0.326258f **FLOATING
C959 a_302_20# 0 0.665072f **FLOATING
C960 a_269_20# 0 0.382299f **FLOATING
C961 a_324_88# 0 0.12884f **FLOATING
C962 b0 0 6.39654f **FLOATING
C963 a0 0 2.56862f **FLOATING
C964 a_810_82# 0 0.382299f **FLOATING
C965 a_734_119# 0 0.665072f **FLOATING
C966 a_769_115# 0 0.100202f **FLOATING
C967 p1 0 6.571078f **FLOATING
C968 a_445_140# 0 0.179875f **FLOATING
C969 a_445_147# 0 0.998982f **FLOATING
C970 pocin 0 0.600283f **FLOATING
C971 a_271_142# 0 0.477455f **FLOATING
C972 a_380_153# 0 0.382299f **FLOATING
C973 a_819_257# 0 0.12884f **FLOATING
C974 a_662_239# 0 0.019534f **FLOATING
C975 a_629_239# 0 0.024435f **FLOATING
C976 a_600_239# 0 0.024435f **FLOATING
C977 a_496_232# 0 0.040245f **FLOATING
C978 cin 0 2.668999f **FLOATING
C979 p0 0 3.844454f **FLOATING
C980 s0 0 0.145867f **FLOATING
C981 a_738_234# 0 0.326258f **FLOATING
C982 a_304_190# 0 0.771781f **FLOATING
C983 a_626_262# 0 0.105692f **FLOATING
C984 a_496_251# 0 0.040245f **FLOATING
C985 p1p0c0 0 0.361176f **FLOATING
C986 a_617_278# 0 0.206277f **FLOATING
C987 a_610_315# 0 0.115609f **FLOATING
C988 a_617_285# 0 1.23327f **FLOATING
C989 a_847_245# 0 0.382299f **FLOATING
C990 a_771_282# 0 0.665072f **FLOATING
C991 a_806_278# 0 0.100202f **FLOATING
C992 a_928_350# 0 0.019534f **FLOATING
C993 a_895_350# 0 0.024435f **FLOATING
C994 a_866_350# 0 0.024435f **FLOATING
C995 a_845_350# 0 0.024435f **FLOATING
C996 a_825_350# 0 0.024435f **FLOATING
C997 a_617_318# 0 0.150155f **FLOATING
C998 a_453_311# 0 1.74716f **FLOATING
C999 a_892_373# 0 0.105692f **FLOATING
C1000 a_271_280# 0 0.477455f **FLOATING
C1001 c4 0 0.15567f **FLOATING
C1002 p3p2p1p0c0 0 0.361176f **FLOATING
C1003 a_776_378# 0 0.019534f **FLOATING
C1004 a_743_378# 0 0.024435f **FLOATING
C1005 a_714_378# 0 0.024435f **FLOATING
C1006 a_693_378# 0 0.024435f **FLOATING
C1007 a_380_291# 0 0.382299f **FLOATING
C1008 a_610_377# 0 0.036687f **FLOATING
C1009 g0 0 10.472128f **FLOATING
C1010 a_304_328# 0 0.771781f **FLOATING
C1011 a_740_401# 0 0.105692f **FLOATING
C1012 a_440_393# 0 0.040245f **FLOATING
C1013 a_610_395# 0 0.040245f **FLOATING
C1014 a_883_389# 0 0.206277f **FLOATING
C1015 a_876_426# 0 0.115609f **FLOATING
C1016 a_883_396# 0 1.73763f **FLOATING
C1017 p2g1 0 0.351373f **FLOATING
C1018 a_610_414# 0 0.040245f **FLOATING
C1019 a_440_412# 0 0.040245f **FLOATING
C1020 a_731_417# 0 0.206277f **FLOATING
C1021 a_724_454# 0 0.115609f **FLOATING
C1022 a_883_429# 0 0.150155f **FLOATING
C1023 p3p2g1 0 0.685912f **FLOATING
C1024 a_731_424# 0 1.49098f **FLOATING
C1025 a_731_457# 0 0.150155f **FLOATING
C1026 p2g1g0 0 0.530242f **FLOATING
C1027 a_883_464# 0 0.148414f **FLOATING
C1028 p3g2 0 0.859094f **FLOATING
C1029 p2p1g0 0 0.15567f **FLOATING
C1030 a_218_418# 0 0.477455f **FLOATING
C1031 a_534_474# 0 2.19469f **FLOATING
C1032 a_397_472# 0 1.74716f **FLOATING
C1033 a_327_429# 0 0.382299f **FLOATING
C1034 a_731_492# 0 0.148414f **FLOATING
C1035 a_884_498# 0 0.144831f **FLOATING
C1036 a_251_466# 0 0.771781f **FLOATING
C1037 a_424_535# 0 0.040245f **FLOATING
C1038 a_594_537# 0 0.040245f **FLOATING
C1039 a_797_547# 0 0.040245f **FLOATING
C1040 a_594_556# 0 0.040245f **FLOATING
C1041 a_424_554# 0 0.040245f **FLOATING
C1042 a_797_566# 0 0.040245f **FLOATING
C1043 a_594_575# 0 0.040245f **FLOATING
C1044 a_797_585# 0 0.040245f **FLOATING
C1045 a_797_604# 0 0.040245f **FLOATING
C1046 a_206_556# 0 0.477455f **FLOATING
C1047 a_315_567# 0 0.382299f **FLOATING
C1048 a_381_614# 0 1.74716f **FLOATING
C1049 a_239_604# 0 0.804448f **FLOATING
C1050 a_518_635# 0 2.19469f **FLOATING
C1051 a_688_664# 0 2.64223f **FLOATING
C1052 w_602_n351# 0 1.34991f **FLOATING
C1053 w_569_n357# 0 1.34991f **FLOATING
C1054 w_401_n374# 0 1.34991f **FLOATING
C1055 w_368_n380# 0 1.34991f **FLOATING
C1056 w_329_n384# 0 1.25349f **FLOATING
C1057 w_292_n385# 0 1.34991f **FLOATING
C1058 w_259_n385# 0 1.34991f **FLOATING
C1059 w_834_n166# 0 1.34991f **FLOATING
C1060 w_801_n166# 0 1.34991f **FLOATING
C1061 w_764_n163# 0 1.25349f **FLOATING
C1062 w_725_n171# 0 1.34991f **FLOATING
C1063 w_692_n177# 0 1.34991f **FLOATING
C1064 w_602_n213# 0 1.34991f **FLOATING
C1065 w_569_n219# 0 1.34991f **FLOATING
C1066 w_401_n240# 0 1.34991f **FLOATING
C1067 w_368_n246# 0 1.34991f **FLOATING
C1068 w_329_n250# 0 1.25349f **FLOATING
C1069 w_292_n251# 0 1.34991f **FLOATING
C1070 w_259_n251# 0 1.34991f **FLOATING
C1071 w_829_n32# 0 1.34991f **FLOATING
C1072 w_796_n32# 0 1.34991f **FLOATING
C1073 w_759_n29# 0 1.25349f **FLOATING
C1074 w_720_n37# 0 1.34991f **FLOATING
C1075 w_687_n43# 0 1.34991f **FLOATING
C1076 w_599_n75# 0 1.34991f **FLOATING
C1077 w_566_n81# 0 1.34991f **FLOATING
C1078 w_400_n106# 0 1.34991f **FLOATING
C1079 w_367_n112# 0 1.34991f **FLOATING
C1080 w_328_n116# 0 1.25349f **FLOATING
C1081 w_291_n117# 0 1.34991f **FLOATING
C1082 w_258_n117# 0 1.34991f **FLOATING
C1083 w_830_114# 0 1.34991f **FLOATING
C1084 w_797_114# 0 1.34991f **FLOATING
C1085 w_760_117# 0 1.25349f **FLOATING
C1086 w_721_109# 0 1.34991f **FLOATING
C1087 w_688_103# 0 1.34991f **FLOATING
C1088 w_602_63# 0 1.34991f **FLOATING
C1089 w_569_57# 0 1.34991f **FLOATING
C1090 w_400_28# 0 1.34991f **FLOATING
C1091 w_367_22# 0 1.34991f **FLOATING
C1092 w_328_18# 0 1.25349f **FLOATING
C1093 w_291_17# 0 1.34991f **FLOATING
C1094 w_258_17# 0 1.34991f **FLOATING
C1095 w_504_133# 0 1.34991f **FLOATING
C1096 w_439_134# 0 1.34991f **FLOATING
C1097 w_439_167# 0 1.34991f **FLOATING
C1098 w_400_185# 0 1.34991f **FLOATING
C1099 w_367_185# 0 1.34991f **FLOATING
C1100 w_291_180# 0 1.34991f **FLOATING
C1101 w_258_174# 0 1.34991f **FLOATING
C1102 w_867_277# 0 1.34991f **FLOATING
C1103 w_834_277# 0 1.34991f **FLOATING
C1104 w_797_280# 0 1.25349f **FLOATING
C1105 w_758_272# 0 1.34991f **FLOATING
C1106 w_725_266# 0 1.34991f **FLOATING
C1107 w_676_271# 0 1.34991f **FLOATING
C1108 w_611_272# 0 1.34991f **FLOATING
C1109 w_611_305# 0 1.34991f **FLOATING
C1110 w_611_340# 0 1.34991f **FLOATING
C1111 w_544_301# 0 1.34991f **FLOATING
C1112 w_506_301# 0 1.34991f **FLOATING
C1113 w_473_301# 0 1.34991f **FLOATING
C1114 w_440_301# 0 1.34991f **FLOATING
C1115 w_400_323# 0 1.34991f **FLOATING
C1116 w_367_323# 0 1.34991f **FLOATING
C1117 w_291_318# 0 1.34991f **FLOATING
C1118 w_258_312# 0 1.34991f **FLOATING
C1119 w_942_382# 0 1.34991f **FLOATING
C1120 w_877_383# 0 1.34991f **FLOATING
C1121 w_877_416# 0 1.34991f **FLOATING
C1122 w_877_451# 0 1.34991f **FLOATING
C1123 w_790_410# 0 1.34991f **FLOATING
C1124 w_725_411# 0 1.34991f **FLOATING
C1125 w_725_444# 0 1.34991f **FLOATING
C1126 w_878_485# 0 1.34991f **FLOATING
C1127 w_725_479# 0 1.34991f **FLOATING
C1128 w_879_518# 0 1.34991f **FLOATING
C1129 w_726_513# 0 1.34991f **FLOATING
C1130 w_658_464# 0 1.34991f **FLOATING
C1131 w_620_464# 0 1.34991f **FLOATING
C1132 w_587_464# 0 1.34991f **FLOATING
C1133 w_554_464# 0 1.34991f **FLOATING
C1134 w_521_464# 0 1.34991f **FLOATING
C1135 w_488_462# 0 1.34991f **FLOATING
C1136 w_450_462# 0 1.34991f **FLOATING
C1137 w_417_462# 0 1.34991f **FLOATING
C1138 w_384_462# 0 1.34991f **FLOATING
C1139 w_347_461# 0 1.34991f **FLOATING
C1140 w_314_461# 0 1.34991f **FLOATING
C1141 w_238_456# 0 1.34991f **FLOATING
C1142 w_205_450# 0 1.34991f **FLOATING
C1143 w_845_654# 0 1.34991f **FLOATING
C1144 w_807_654# 0 1.34991f **FLOATING
C1145 w_774_654# 0 1.34991f **FLOATING
C1146 w_741_654# 0 1.34991f **FLOATING
C1147 w_708_654# 0 1.34991f **FLOATING
C1148 w_675_654# 0 1.34991f **FLOATING
C1149 w_642_625# 0 1.34991f **FLOATING
C1150 w_604_625# 0 1.34991f **FLOATING
C1151 w_571_625# 0 1.34991f **FLOATING
C1152 w_538_625# 0 1.34991f **FLOATING
C1153 w_505_625# 0 1.34991f **FLOATING
C1154 w_472_604# 0 1.34991f **FLOATING
C1155 w_434_604# 0 1.34991f **FLOATING
C1156 w_401_604# 0 1.34991f **FLOATING
C1157 w_368_604# 0 1.34991f **FLOATING
C1158 w_335_599# 0 1.34991f **FLOATING
C1159 w_302_599# 0 1.34991f **FLOATING
C1160 w_226_594# 0 1.34991f **FLOATING
C1161 w_193_588# 0 1.34991f **FLOATING
