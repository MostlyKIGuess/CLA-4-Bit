* OR Testing Code
* TSMC 180nm Technology Parameters
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Supply
Vdd vdd gnd 'SUPPLY'

* Test Signals
Vclk b gnd PULSE(0 'SUPPLY' 0 0.001n 0.01n 10n 20n)
Vd a gnd PULSE(0 'SUPPLY' 0n 0.001n 0.01n 35n 70n)



* OR Gate Subcircuit
.subckt or a b y vdd gnd
    * NOR
    Mn1 ybar a gnd gnd CMOSN L={2*LAMBDA} W={width_N} AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Mn2 ybar b gnd gnd CMOSN L={2*LAMBDA} W={width_N} AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Mp1 ybar b c vdd CMOSP L={2*LAMBDA} W={width_P} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    Mp2 c a vdd vdd CMOSP L={2*LAMBDA} W={width_P} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    * inverter
    Mn4 y ybar gnd gnd CMOSN L={2*LAMBDA} W={width_N} AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Mp3 y ybar vdd vdd CMOSP L={2*LAMBDA} W={width_P} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends or
* Instantiate the OR Gate
Xor1 a b out vdd gnd or

.control
  set hcopypscolor = 1
  set color0 = white
  set color1 = black
  set color2 = red
  set color3 = blue
  set color4 = brown
  set color5 = magenta
  set color6 = cyan
  set color7 = green
  tran 1n 200n
    plot a 2+b 4+out
.endc


