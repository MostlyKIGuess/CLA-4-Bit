* SPICE3 file created from or.ext - technology: scmos

.option scale=1u

M1000 ybar b gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 ybar c gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 ybar c a_n75_7# w_n81_1# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1003 y ybar vdd w_n16_0# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 vdd b a_n75_7# w_n81_34# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1005 y ybar gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
C0 w_n81_34# vdd 1.41f
C1 gnd ybar 0.808f
C2 w_n81_1# a_n75_7# 2.444f
C3 w_n16_0# vdd 1.128f
C4 c w_n81_1# 2.312f
C5 ybar w_n16_0# 1.014f
C6 w_n81_34# a_n75_7# 1.128f
C7 w_n16_0# y 1.88f
C8 w_n81_34# b 1.482f
C9 w_n81_1# ybar 1.88f
C10 gnd 0 11.561999f **FLOATING
C11 y 0 4.324f **FLOATING
C12 c 0 8.299999f **FLOATING
C13 a_n75_7# 0 4.888f **FLOATING
C14 b 0 24.082f **FLOATING
C15 ybar 0 19.995f **FLOATING
C16 vdd 0 13.536f **FLOATING
