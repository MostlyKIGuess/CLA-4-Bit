* NGSPICE file created from testing.ext - technology: scmos

.option scale=1u

M1000 a_445_147# g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 a_691_n240# a_615_n203# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_615_n203# a_582_n251# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 p2g1 a_327_429# vdd w_347_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_594_575# p1 a_594_556# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1005 a_440_412# p1 a_440_393# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 p1p0c0 a_453_311# vdd w_544_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 a3 a_338_n335# a_303_n382# w_329_n384# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 a_848_2# p2 c2 w_835_n8# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1009 a_518_635# p3 vdd w_505_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_731_457# p2p1p0c0 a_731_417# w_725_444# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1011 b2 a2 a_303_n248# w_368_n246# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1012 gnd a_303_n248# a_270_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 p3p2g1 a_381_614# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 p2p1p0c0 a_534_474# vdd w_658_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 a_610_395# p1 a_610_377# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1016 gnd a_325_n180# a_303_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1017 a_815_n46# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1018 a_518_635# g0 a_594_575# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_940_n169# a_864_n132# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1020 s2 a_924_n35# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1021 vdd a0 a_345_92# w_400_28# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 vdd a_302_20# a_269_20# w_291_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a_346_n176# b2 a_303_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1024 g0 a_691_36# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1025 a_825_350# p3p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1026 a_847_245# a_771_282# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 a_304_190# a_271_142# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1028 a_884_498# p3g2 a_883_464# w_878_485# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1029 g3 a_691_n378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 a_731_492# p2p1g0 a_731_457# w_725_479# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 a_831_148# a_879_123# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 a_615_n341# a3 b3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1033 a_831_148# a_866_144# p1 w_857_146# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1034 a_798_100# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1035 a_315_567# a_239_604# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 g2 a_691_n240# vdd w_711_n208# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1037 a_582_n251# a2 vdd w_569_n219# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1038 p3g2 a_315_567# vdd w_335_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1039 vdd g3 a_884_498# w_879_518# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 a_825_350# p3p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1041 pocin a_380_153# vdd w_400_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1042 vdd a_269_20# p0 w_258_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1043 a_218_418# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 a_380_153# a_304_190# vdd w_367_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 b1 a1 a_302_n114# w_367_n112# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 a_691_36# a_615_73# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1047 a_825_350# p3p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 a_271_280# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1049 a_907_111# a_831_148# vdd w_894_143# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 s2 a_924_n35# vdd w_944_n3# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1051 p3p2p1g0 a_518_635# vdd w_642_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 a_615_n203# a_582_n251# b2 w_602_n213# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_239_604# a_206_556# g2 w_226_594# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1054 a_304_190# a_271_142# cin w_291_180# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1055 a_612_n65# a_579_n113# b1 w_599_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_582_25# a0 vdd w_569_57# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 p2p1g0 a_397_472# vdd w_488_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 c3 a_693_378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 a_440_393# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1060 a_612_n65# a_579_n113# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1061 a_924_n35# a_848_2# vdd w_911_n3# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_688_664# p0 vdd w_774_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 a_445_147# pocin gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1064 p2g1 a_327_429# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 a_600_239# p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 s3 a_940_n169# vdd w_960_n137# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1067 a_327_429# a_251_466# vdd w_314_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_848_2# a_896_n23# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1069 a_688_664# cin vdd w_807_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 a_693_378# p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1071 a_251_466# p2 g1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_346_n310# b3 a_303_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 a_688_n102# a_612_n65# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_738_234# p0 vdd w_725_266# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_924_n35# a_848_2# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 p3p2g1 a_381_614# vdd w_472_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1077 a_206_556# p3 vdd w_193_588# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1078 a_424_535# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1079 g2 a_691_n240# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1080 a_610_377# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1081 s0 a_847_245# vdd w_867_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_582_n389# a3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1083 a_691_n378# a_615_n341# vdd w_678_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1084 a_864_n132# a_912_n157# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1085 vdd a2 a_346_n176# w_401_n240# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_615_n203# a2 b2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1087 g1 a_688_n102# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1088 c4 a_825_350# vdd w_942_382# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_424_554# p2 a_424_535# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 a_453_311# p0 vdd w_473_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_831_n180# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_315_567# a_239_604# vdd w_302_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 p3p2p1p0c0 a_688_664# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1094 a_771_282# p0 cin w_758_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 a_271_142# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_612_n65# a1 b1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1097 a_534_474# cin vdd w_620_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_534_474# p0 vdd w_587_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1099 a_453_311# cin vdd w_506_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_271_280# p1 vdd w_258_312# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_693_378# p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1102 a_381_614# g1 a_424_554# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_883_429# p3p2p1g0 a_883_389# w_877_416# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 c1 a_445_147# vdd w_504_133# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_304_328# a_271_280# g0 w_291_318# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_825_350# p3g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 a_688_664# p1 vdd w_741_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_797_604# p0 a_797_585# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 vdd a_269_n114# p1 w_258_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1110 p1g0 a_380_291# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 a_345_n42# b1 a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_327_429# a_251_466# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1113 a1 a_337_n67# a_302_n114# w_328_n116# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 s1 a_907_111# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1115 a_693_378# p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_380_291# a_304_328# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 c2 a_600_239# vdd w_676_271# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1118 gnd a_324_88# a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 b3 a3 a_303_n382# w_368_n380# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1120 a_688_n102# a_612_n65# vdd w_675_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 gnd a_324_n46# a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1122 a_815_n46# p2 vdd w_802_n14# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 vdd a3 a_346_n310# w_401_n374# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1124 a_615_73# a_582_25# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 p1p0c0 a_453_311# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1126 a_345_92# b0 a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 a_688_664# cin a_797_604# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1128 vdd g2 a_731_492# w_726_513# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1129 a_883_464# p3p2g1 a_883_429# w_877_451# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 a_693_378# g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1131 g1 a_688_n102# vdd w_708_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_831_148# c1 a_798_100# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_864_n132# p3 c3 w_851_n142# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1134 a_304_328# p1 g0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1135 a_771_282# a_819_257# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1136 a_518_635# p1 vdd w_571_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1137 a_397_472# g0 vdd w_450_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1138 a_579_n113# a1 vdd w_566_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_797_547# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_496_251# p0 a_496_232# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_848_2# a_883_n2# p2 w_874_0# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 g0 a_691_36# vdd w_711_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_847_245# a_771_282# vdd w_834_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1147 vdd a_270_n248# p2 w_259_n251# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1148 a_579_n113# a1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1149 a_239_604# a_206_556# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1150 a_797_566# p2 a_797_547# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 a_453_311# cin a_496_251# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1152 a_453_311# p1 vdd w_440_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_798_100# p1 vdd w_785_132# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1154 gnd a3 a_346_n310# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1155 a_534_474# p1 vdd w_554_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 a_304_328# a_271_280# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_445_147# g0 a_445_140# w_439_134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1158 a_940_n169# a_864_n132# vdd w_927_n137# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1159 a_797_585# p1 a_797_566# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1160 a_864_n132# c3 a_831_n180# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1161 gnd a_302_n114# a_269_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_691_36# a_615_73# vdd w_678_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1163 s3 a_940_n169# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_864_n132# a_899_n136# p3 w_890_n134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1165 gnd a_269_n114# p1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1166 a_381_614# g1 vdd w_434_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1167 vdd a_303_n248# a_270_n248# w_292_n251# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 pocin a_380_153# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 a_848_2# c2 a_815_n46# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1170 a_380_153# a_304_190# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 a_831_148# p1 c1 w_818_138# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1172 a_688_664# p3 vdd w_675_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 g3 a_691_n378# vdd w_711_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_907_111# a_831_148# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1175 p1g0 a_380_291# vdd w_400_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1176 c2 a_600_239# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 a_615_73# a0 b0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1178 a0 a_337_67# a_302_20# w_328_18# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_380_291# a_304_328# vdd w_367_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1180 vdd a_270_n382# p3 w_259_n385# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1181 a_582_25# a0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1182 a_688_664# p2 vdd w_708_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 p2p1g0 a_397_472# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1184 gnd a2 a_346_n176# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1185 vdd pocin a_445_140# w_439_167# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 c3 a_693_378# vdd w_790_410# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1187 a_304_190# p0 cin Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_251_466# a_218_418# g1 w_238_456# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 vdd a1 a_345_n42# w_400_n106# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# g0 a_440_412# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 a_691_n378# a_615_n341# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1192 a_615_n341# a_582_n389# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1193 a_397_472# p2 vdd w_384_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 vdd a_303_n382# a_270_n382# w_292_n385# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1195 vdd a_302_n114# a_269_n114# w_291_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_617_318# p1g0 a_617_278# w_611_305# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 a_771_282# a_806_278# p0 w_797_280# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_738_234# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1199 a_691_n240# a_615_n203# vdd w_678_n208# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_518_635# p2 vdd w_538_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1201 a_496_232# p1 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 b0 a0 a_302_20# w_367_22# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_397_472# p1 vdd w_417_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_206_556# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1205 gnd a_270_n382# p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 a_610_414# p0 a_610_395# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 p3p2p1p0c0 a_688_664# vdd w_845_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1208 a_271_142# p0 vdd w_258_174# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1209 a_582_n251# a2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 a_534_474# p2 vdd w_521_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1211 s0 a_847_245# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1212 vdd g1 a_617_318# w_611_340# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 c4 a_825_350# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 gnd a0 a_345_92# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1215 gnd a1 a_345_n42# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 gnd a_302_20# a_269_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1217 a_381_614# p2 vdd w_401_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1218 a_534_474# cin a_610_414# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1219 a2 a_338_n201# a_303_n248# w_329_n250# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1220 a_251_466# a_218_418# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1221 a_771_282# cin a_738_234# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1222 a_381_614# p3 vdd w_368_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1223 p3g2 a_315_567# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1224 a_594_537# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1225 a_600_239# g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1226 a_615_73# a_582_25# b0 w_602_63# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1227 a_582_n389# a3 vdd w_569_n357# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1228 a_239_604# p3 g2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1229 gnd a_325_n314# a_303_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1230 gnd a_303_n382# a_270_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1231 a_218_418# p2 vdd w_205_450# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1232 a_825_350# g3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1233 a_600_239# p1p0c0 a_617_278# w_611_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1234 s1 a_907_111# vdd w_927_143# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1235 c1 a_445_147# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1236 p3p2p1g0 a_518_635# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1237 a_693_378# p2g1 a_731_417# w_725_411# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1238 a_831_n180# p3 vdd w_818_n148# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1239 a_600_239# p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1240 gnd a_270_n248# p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1241 a_594_556# p2 a_594_537# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1242 gnd a_269_20# p0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1243 a_615_n341# a_582_n389# b3 w_602_n351# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 w_658_464# vdd 1.128f
C1 a_825_350# gnd 3.232f
C2 w_440_301# a_453_311# 2.45f
C3 w_368_n246# b2 1.88f
C4 w_292_n251# a_270_n248# 1.88f
C5 w_911_n3# vdd 1.128f
C6 w_620_464# vdd 1.128f
C7 w_401_604# p2 1.014f
C8 w_259_n251# a_270_n248# 1.014f
C9 w_678_n208# a_615_n203# 1.014f
C10 p3 vdd 2.52f
C11 w_587_464# vdd 1.128f
C12 w_417_462# p1 1.014f
C13 w_620_464# cin 1.014f
C14 w_602_n213# a_615_n203# 2.82f
C15 w_569_n219# a2 1.014f
C16 w_554_464# vdd 1.128f
C17 w_401_n240# a2 1.014f
C18 w_802_n14# vdd 1.128f
C19 g0 p1p0c0 0.18f
C20 w_259_n385# p3 1.88f
C21 w_818_138# c1 1.88f
C22 w_521_464# vdd 1.128f
C23 w_291_318# a_271_280# 1.014f
C24 w_587_464# p0 1.014f
C25 w_711_68# vdd 1.128f
C26 w_368_n246# a2 1.17f
C27 w_488_462# vdd 1.128f
C28 w_400_323# a_380_291# 1.014f
C29 w_258_312# a_271_280# 1.88f
C30 g0 p1g0 1.01f
C31 w_678_68# vdd 1.128f
C32 w_960_n137# s3 1.88f
C33 w_329_n250# a2 1.128f
C34 w_226_594# g2 2.268f
C35 w_845_654# a_688_664# 1.014f
C36 w_504_133# c1 1.88f
C37 w_927_143# a_907_111# 1.014f
C38 w_785_132# a_798_100# 1.88f
C39 w_708_n70# g1 1.88f
C40 c3 a_912_n157# 0.54f
C41 w_450_462# vdd 1.128f
C42 w_367_323# a_380_291# 1.88f
C43 w_193_588# g2 1.064f
C44 w_807_654# a_688_664# 3.59f
C45 w_894_143# a_907_111# 1.88f
C46 w_417_462# vdd 1.128f
C47 w_400_323# g0 1.33f
C48 w_942_382# c4 1.88f
C49 w_569_57# vdd 1.128f
C50 w_774_654# a_688_664# 3.59f
C51 a_206_556# g2 0.846f
C52 w_894_143# a_831_148# 1.014f
C53 b2 a_346_n176# 1.08f
C54 w_384_462# vdd 1.128f
C55 a_693_378# gnd 2.424f
C56 w_367_323# g0 1.33f
C57 w_400_28# vdd 1.128f
C58 w_741_654# a_688_664# 3.59f
C59 w_857_146# a_831_148# 1.128f
C60 b2 a_303_n248# 6.03f
C61 w_347_461# vdd 1.128f
C62 b0 a_345_92# 1.08f
C63 w_877_383# p3p2p1p0c0 2.202f
C64 w_367_323# a_304_328# 1.014f
C65 w_291_318# g0 1.128f
C66 a_381_614# p2 0.19f
C67 w_851_n142# c3 1.88f
C68 w_708_654# a_688_664# 3.59f
C69 w_439_134# a_445_140# 2.444f
C70 w_504_133# a_445_147# 1.014f
C71 w_818_138# a_831_148# 2.162f
C72 w_857_146# a_866_144# 1.17f
C73 w_314_461# vdd 1.128f
C74 c1 a_879_123# 0.54f
C75 b0 a_302_20# 6.03f
C76 w_291_318# a_304_328# 2.82f
C77 w_960_n137# a_940_n169# 1.014f
C78 w_675_654# a_688_664# 2.45f
C79 w_642_625# a_518_635# 1.014f
C80 w_439_134# a_445_147# 1.88f
C81 w_439_167# a_445_140# 1.128f
C82 w_857_146# p1 1.128f
C83 a_239_604# g2 0.786f
C84 b2 a_325_n180# 0.54f
C85 w_741_654# p1 1.014f
C86 a_534_474# p1 0.19f
C87 w_927_n137# a_940_n169# 1.88f
C88 a_518_635# p2 0.19f
C89 w_291_17# vdd 1.128f
C90 w_818_n148# a_831_n180# 1.88f
C91 w_604_625# a_518_635# 3.59f
C92 w_818_138# p1 1.17f
C93 b1 gnd 2.314f
C94 w_205_450# vdd 1.128f
C95 b0 a_324_88# 0.54f
C96 a_688_664# p2 0.19f
C97 w_258_17# vdd 1.128f
C98 a_397_472# p1 0.19f
C99 w_927_n137# a_864_n132# 1.014f
C100 w_571_625# a_518_635# 3.59f
C101 w_785_132# p1 1.014f
C102 w_845_654# vdd 1.128f
C103 g1 a_615_n203# 2.97f
C104 w_890_n134# a_864_n132# 1.128f
C105 w_927_143# vdd 1.128f
C106 w_472_604# a_381_614# 1.014f
C107 w_538_625# a_518_635# 3.59f
C108 b1 vdd 0.9f
C109 w_807_654# vdd 1.128f
C110 w_790_410# c3 1.88f
C111 a0 b0 4.458f
C112 w_894_143# vdd 1.128f
C113 w_851_n142# a_864_n132# 2.162f
C114 w_890_n134# a_899_n136# 1.17f
C115 w_434_604# a_381_614# 3.59f
C116 w_258_17# p0 1.88f
C117 w_505_625# a_518_635# 2.45f
C118 a1 vdd 2.52f
C119 w_676_271# c2 1.88f
C120 w_774_654# vdd 1.128f
C121 w_890_n134# p3 1.128f
C122 w_807_654# cin 1.014f
C123 w_401_604# a_381_614# 3.59f
C124 a2 b2 3.468f
C125 a_612_n65# vdd 1.35f
C126 w_741_654# vdd 1.128f
C127 w_877_383# a_883_389# 2.444f
C128 w_571_625# p1 1.014f
C129 w_851_n142# p3 1.17f
C130 g0 a_380_291# 1.01f
C131 w_439_167# pocin 1.482f
C132 w_368_604# a_381_614# 2.45f
C133 w_335_599# a_315_567# 1.014f
C134 a_615_n203# b2 1.91f
C135 w_708_654# vdd 1.128f
C136 g1 p3 83.43f
C137 w_818_n148# p3 1.014f
C138 w_774_654# p0 1.014f
C139 a_534_474# cin 0.19f
C140 w_877_416# a_883_389# 1.128f
C141 w_942_382# a_825_350# 1.014f
C142 w_785_132# vdd 1.128f
C143 w_302_599# a_315_567# 1.88f
C144 w_226_594# a_206_556# 1.014f
C145 w_400_185# pocin 1.88f
C146 a_615_73# b0 1.91f
C147 w_675_654# vdd 1.128f
C148 g2 gnd 30.06f
C149 w_877_383# a_825_350# 1.88f
C150 w_877_416# p3p2p1g0 1.482f
C151 w_504_133# vdd 1.128f
C152 w_834_277# vdd 1.128f
C153 a_534_474# p0 0.19f
C154 w_193_588# a_206_556# 1.88f
C155 w_642_625# vdd 1.128f
C156 a_304_328# g0 1.35f
C157 w_302_599# a_239_604# 1.014f
C158 w_400_185# a_380_153# 1.014f
C159 p2 vdd 2.52f
C160 g2 vdd 2.068f
C161 w_604_625# vdd 1.128f
C162 w_439_167# vdd 1.41f
C163 w_367_185# a_380_153# 1.88f
C164 w_291_180# a_271_142# 1.014f
C165 w_226_594# a_239_604# 2.82f
C166 a_864_n132# c3 6.03f
C167 w_571_625# vdd 1.128f
C168 w_400_185# vdd 1.128f
C169 w_258_174# a_271_142# 1.88f
C170 a_251_466# vdd 1.89f
C171 w_538_625# vdd 1.128f
C172 w_367_185# vdd 1.128f
C173 w_708_n70# a_688_n102# 1.014f
C174 w_711_n208# g2 1.88f
C175 w_505_625# vdd 1.128f
C176 w_725_411# p2g1 2.202f
C177 w_675_n70# a_688_n102# 1.88f
C178 w_599_n75# a_579_n113# 1.014f
C179 w_472_604# vdd 1.128f
C180 w_566_n81# a_579_n113# 1.88f
C181 w_258_174# vdd 1.128f
C182 w_291_180# cin 1.128f
C183 w_434_604# vdd 1.128f
C184 a_831_148# c1 6.03f
C185 w_867_277# vdd 1.128f
C186 w_877_416# a_883_429# 1.41f
C187 w_401_604# vdd 1.128f
C188 w_238_456# g1 2.724f
C189 w_877_451# a_883_429# 1.41f
C190 w_725_411# a_731_417# 2.444f
C191 w_328_n116# a_337_n67# 1.17f
C192 w_258_174# p0 1.014f
C193 w_711_68# g0 1.88f
C194 b0 gnd 1.91f
C195 w_368_604# vdd 1.128f
C196 w_205_450# g1 1.596f
C197 w_400_n106# a_345_n42# 1.88f
C198 w_725_444# a_731_417# 1.128f
C199 w_877_451# p3p2g1 1.482f
C200 w_367_185# a_304_190# 1.014f
C201 w_335_599# vdd 1.128f
C202 w_725_444# p2p1p0c0 1.482f
C203 w_450_462# g0 1.014f
C204 w_291_180# a_304_190# 2.82f
C205 w_867_277# s0 1.88f
C206 b0 vdd 0.9f
C207 w_302_599# vdd 1.128f
C208 w_790_410# a_693_378# 1.014f
C209 w_367_n112# a_302_n114# 2.162f
C210 w_834_277# a_847_245# 1.88f
C211 a0 vdd 2.52f
C212 g1 a1 16.199999f
C213 g2 a_615_n341# 1.485f
C214 w_725_411# a_693_378# 1.88f
C215 w_259_n251# p2 1.88f
C216 w_328_n116# a_302_n114# 1.128f
C217 a_218_418# g1 1.212f
C218 w_834_277# a_771_282# 1.014f
C219 w_193_588# vdd 1.128f
C220 w_877_451# a_883_464# 1.598f
C221 w_291_n117# a_302_n114# 1.014f
C222 a_518_635# p1 0.19f
C223 w_725_444# a_731_457# 1.41f
C224 w_845_654# p3p2p1p0c0 1.88f
C225 w_291_n117# a_269_n114# 1.88f
C226 w_599_n75# b1 1.128f
C227 a_688_664# p1 0.19f
C228 w_658_464# p2p1p0c0 1.88f
C229 w_258_n117# a_269_n114# 1.014f
C230 w_675_n70# a_612_n65# 1.014f
C231 a_615_73# vdd 1.35f
C232 a_445_147# gnd 0.808f
C233 w_725_479# a_731_457# 1.41f
C234 w_400_n106# b1 1.71f
C235 w_599_n75# a_612_n65# 2.82f
C236 w_566_n81# a1 1.014f
C237 g1 p2 3.825f
C238 a_239_604# vdd 1.89f
C239 w_878_485# a_883_464# 1.41f
C240 w_725_479# p2p1g0 1.482f
C241 w_367_n112# b1 1.88f
C242 w_400_n106# a1 1.014f
C243 w_878_485# p3g2 1.482f
C244 w_944_n3# s2 1.88f
C245 w_367_n112# a1 1.17f
C246 w_867_277# a_847_245# 1.014f
C247 w_711_n346# g3 1.88f
C248 a_251_466# g1 1.212f
C249 w_328_n116# a1 1.128f
C250 w_711_n346# vdd 1.128f
C251 w_347_461# p2g1 1.88f
C252 a_688_664# cin 0.19f
C253 w_678_n346# vdd 1.128f
C254 a_688_664# p0 0.19f
C255 a_397_472# g0 0.19f
C256 p1 vdd 2.52f
C257 w_434_604# g1 1.014f
C258 w_835_n8# c2 1.88f
C259 w_504_133# g0 1.33f
C260 c2 a_896_n23# 0.54f
C261 w_711_n346# a_691_n378# 1.014f
C262 w_569_n357# vdd 1.128f
C263 w_439_134# g0 2.943f
C264 w_678_n346# a_691_n378# 1.88f
C265 w_401_n374# vdd 1.128f
C266 w_602_n351# a_582_n389# 1.014f
C267 w_604_625# g0 1.014f
C268 w_725_479# a_731_492# 1.598f
C269 w_658_464# a_534_474# 1.014f
C270 w_802_n14# a_815_n46# 1.88f
C271 w_944_n3# a_924_n35# 1.014f
C272 w_569_n357# a_582_n389# 1.88f
C273 w_620_464# a_534_474# 3.59f
C274 w_878_485# a_884_498# 1.598f
C275 w_488_462# p2p1g0 1.88f
C276 w_911_n3# a_924_n35# 1.88f
C277 w_587_464# a_534_474# 3.59f
C278 w_726_513# a_731_492# 1.41f
C279 w_911_n3# a_848_2# 1.014f
C280 w_292_n385# vdd 1.128f
C281 w_329_n384# a_338_n335# 1.17f
C282 cin a_819_257# 0.54f
C283 w_879_518# a_884_498# 1.41f
C284 w_726_513# g2 1.482f
C285 w_554_464# a_534_474# 3.59f
C286 w_874_0# a_848_2# 1.128f
C287 cin vdd 1.26f
C288 w_675_654# p3 1.014f
C289 w_259_n385# vdd 1.128f
C290 w_401_n374# a_346_n310# 1.88f
C291 w_521_464# a_534_474# 2.45f
C292 w_642_625# p3p2p1g0 1.88f
C293 w_835_n8# a_848_2# 2.162f
C294 w_874_0# a_883_n2# 1.17f
C295 w_725_266# vdd 1.128f
C296 p0 vdd 2.52f
C297 b1 a_345_n42# 1.08f
C298 w_758_272# cin 1.88f
C299 w_797_280# p0 1.128f
C300 w_711_n208# vdd 1.128f
C301 w_874_0# p2 1.128f
C302 w_676_271# vdd 1.128f
C303 b1 a_302_n114# 6.03f
C304 w_758_272# p0 1.17f
C305 w_368_n380# a_303_n382# 2.162f
C306 w_678_n208# vdd 1.128f
C307 g2 p3 1.575f
C308 w_602_n351# b3 1.128f
C309 w_488_462# a_397_472# 1.014f
C310 w_835_n8# p2 1.17f
C311 w_725_266# p0 1.014f
C312 w_678_n346# a_615_n341# 1.014f
C313 w_329_n384# a_303_n382# 1.128f
C314 w_450_462# a_397_472# 3.59f
C315 w_802_n14# p2 1.014f
C316 a_381_614# g1 0.19f
C317 b1 a_324_n46# 0.54f
C318 a_304_190# vdd 1.89f
C319 w_440_301# p1 1.014f
C320 w_521_464# p2 1.014f
C321 w_401_n374# b3 1.71f
C322 w_602_n351# a_615_n341# 2.82f
C323 w_569_n357# a3 1.014f
C324 w_292_n385# a_303_n382# 1.014f
C325 w_569_n219# vdd 1.128f
C326 w_417_462# a_397_472# 3.59f
C327 b3 gnd 1.73f
C328 w_611_340# vdd 1.88f
C329 w_401_n240# vdd 1.128f
C330 w_368_n380# b3 1.88f
C331 w_292_n385# a_270_n382# 1.88f
C332 w_401_n374# a3 1.014f
C333 w_505_625# p3 1.014f
C334 w_725_266# a_738_234# 1.88f
C335 w_384_462# a_397_472# 2.45f
C336 w_544_301# vdd 1.128f
C337 w_368_n380# a3 1.17f
C338 w_259_n385# a_270_n382# 1.014f
C339 w_238_456# a_218_418# 1.014f
C340 b3 vdd 0.72f
C341 w_506_301# vdd 1.128f
C342 a_600_239# gnd 1.616f
C343 w_329_n384# a3 1.128f
C344 w_347_461# a_327_429# 1.014f
C345 w_205_450# a_218_418# 1.88f
C346 a3 vdd 2.52f
C347 w_473_301# vdd 1.128f
C348 w_258_312# p1 1.014f
C349 w_506_301# cin 1.014f
C350 w_384_462# p2 1.014f
C351 g0 c1 1.01f
C352 w_292_n251# vdd 1.128f
C353 w_602_63# a_582_25# 1.014f
C354 w_711_68# a_691_36# 1.014f
C355 w_314_461# a_327_429# 1.88f
C356 a_615_n341# vdd 1.08f
C357 w_440_301# vdd 1.128f
C358 a1 b1 4.008f
C359 w_259_n251# vdd 1.128f
C360 w_368_604# p3 1.014f
C361 w_678_68# a_691_36# 1.88f
C362 w_569_57# a_582_25# 1.88f
C363 w_400_323# vdd 1.128f
C364 a_848_2# c2 6.03f
C365 a_612_n65# b1 2.674f
C366 w_611_272# p1p0c0 2.202f
C367 w_473_301# p0 1.014f
C368 w_960_n137# vdd 1.128f
C369 b3 a_346_n310# 1.08f
C370 w_367_323# vdd 1.128f
C371 w_797_280# a_771_282# 1.128f
C372 w_611_272# a_617_278# 2.444f
C373 w_927_n137# vdd 1.128f
C374 w_328_18# a_337_67# 1.17f
C375 b3 a_303_n382# 6.03f
C376 g1 gnd 15.03f
C377 w_758_272# a_771_282# 2.162f
C378 w_611_305# a_617_278# 1.128f
C379 w_676_271# a_600_239# 1.014f
C380 w_797_280# a_806_278# 1.17f
C381 w_205_450# p2 1.014f
C382 g0 a_445_147# 0.72f
C383 a_771_282# cin 6.03f
C384 a_518_635# g0 0.19f
C385 w_314_461# a_251_466# 1.014f
C386 w_258_312# vdd 1.128f
C387 w_544_301# p1p0c0 1.88f
C388 w_193_588# p3 1.014f
C389 w_611_272# a_600_239# 1.88f
C390 w_611_305# p1g0 1.482f
C391 w_472_604# p3p2g1 1.88f
C392 w_238_456# a_251_466# 2.82f
C393 w_400_28# a_345_92# 1.88f
C394 b3 a_325_n314# 0.54f
C395 g1 vdd 2.472f
C396 w_942_382# vdd 1.128f
C397 w_818_n148# vdd 1.128f
C398 w_708_n70# vdd 1.128f
C399 w_711_n208# a_691_n240# 1.014f
C400 w_602_63# b0 1.128f
C401 w_367_22# a_302_20# 2.162f
C402 a3 b3 3.738f
C403 b2 gnd 1.91f
C404 w_678_n208# a_691_n240# 1.88f
C405 w_602_n213# a_582_n251# 1.014f
C406 a_453_311# cin 0.19f
C407 w_675_n70# vdd 1.128f
C408 w_328_18# a_302_20# 1.128f
C409 a_615_n341# b3 1.91f
C410 w_569_n219# a_582_n251# 1.88f
C411 a_453_311# p0 0.19f
C412 w_708_654# p2 1.014f
C413 w_400_28# b0 1.71f
C414 w_291_17# a_302_20# 1.014f
C415 w_569_57# a0 1.014f
C416 b2 vdd 0.9f
C417 w_790_410# vdd 1.128f
C418 w_611_305# a_617_318# 1.41f
C419 w_566_n81# vdd 1.128f
C420 w_367_22# b0 1.88f
C421 w_291_17# a_269_20# 1.88f
C422 w_400_28# a0 1.014f
C423 w_258_n117# p1 1.88f
C424 w_611_340# a_617_318# 1.41f
C425 w_400_323# p1g0 1.88f
C426 w_329_n250# a_338_n201# 1.17f
C427 w_400_n106# vdd 1.128f
C428 w_367_22# a0 1.17f
C429 w_258_17# a_269_20# 1.014f
C430 w_678_68# a_615_73# 1.014f
C431 w_611_340# g1 1.482f
C432 w_401_n240# a_346_n176# 1.88f
C433 w_328_18# a0 1.128f
C434 w_602_63# a_615_73# 2.82f
C435 g0 vdd 4.29f
C436 a2 vdd 2.52f
C437 w_879_518# g3 1.482f
C438 a_304_328# vdd 1.89f
C439 w_538_625# p2 1.014f
C440 w_544_301# a_453_311# 1.014f
C441 w_291_n117# vdd 1.128f
C442 w_602_n213# b2 1.128f
C443 w_368_n246# a_303_n248# 2.162f
C444 w_335_599# p3g2 1.88f
C445 a_615_n203# vdd 1.35f
C446 w_879_518# vdd 1.88f
C447 w_554_464# p1 1.014f
C448 w_506_301# a_453_311# 3.59f
C449 w_258_n117# vdd 1.128f
C450 w_329_n250# a_303_n248# 1.128f
C451 w_726_513# vdd 1.88f
C452 w_473_301# a_453_311# 3.59f
C453 w_401_n240# b2 1.71f
C454 w_292_n251# a_303_n248# 1.014f
C455 w_944_n3# vdd 1.128f
C456 w_927_143# s1 1.88f
C457 gnd 0 1.292547p $ **FLOATING
C458 g3 0 65.881004f $ **FLOATING
C459 vdd 0 0.952454p $ **FLOATING
C460 a_338_n335# 0 3.508f $ **FLOATING
C461 a_582_n389# 0 18.082f $ **FLOATING
C462 a_691_n378# 0 14.266f $ **FLOATING
C463 a_346_n310# 0 14.946f $ **FLOATING
C464 a_303_n382# 0 31.139002f $ **FLOATING
C465 a_270_n382# 0 14.266f $ **FLOATING
C466 a_325_n314# 0 4.916f $ **FLOATING
C467 b3 0 85.516f $ **FLOATING
C468 a3 0 0.140213p $ **FLOATING
C469 a_615_n341# 0 44.863f $ **FLOATING
C470 a_912_n157# 0 4.916f $ **FLOATING
C471 a_338_n201# 0 3.508f $ **FLOATING
C472 a_582_n251# 0 18.082f $ **FLOATING
C473 a_691_n240# 0 14.266f $ **FLOATING
C474 a_346_n176# 0 14.946f $ **FLOATING
C475 a_303_n248# 0 31.139002f $ **FLOATING
C476 a_270_n248# 0 14.266f $ **FLOATING
C477 a_325_n180# 0 4.916f $ **FLOATING
C478 b2 0 85.212006f $ **FLOATING
C479 s3 0 3.76f $ **FLOATING
C480 c3 0 17.83f $ **FLOATING
C481 a_831_n180# 0 14.946f $ **FLOATING
C482 a2 0 0.137957p $ **FLOATING
C483 a_615_n203# 0 44.863f $ **FLOATING
C484 a_940_n169# 0 14.266f $ **FLOATING
C485 a_864_n132# 0 31.139002f $ **FLOATING
C486 a_899_n136# 0 3.508f $ **FLOATING
C487 p3 0 0.378435p $ **FLOATING
C488 a_896_n23# 0 4.916f $ **FLOATING
C489 a_337_n67# 0 3.508f $ **FLOATING
C490 a_579_n113# 0 18.082f $ **FLOATING
C491 a_688_n102# 0 14.266f $ **FLOATING
C492 a_345_n42# 0 14.946f $ **FLOATING
C493 a_302_n114# 0 31.139002f $ **FLOATING
C494 a_269_n114# 0 14.266f $ **FLOATING
C495 a_324_n46# 0 4.916f $ **FLOATING
C496 s2 0 3.76f $ **FLOATING
C497 c2 0 17.83f $ **FLOATING
C498 a_815_n46# 0 14.946f $ **FLOATING
C499 b1 0 88.200005f $ **FLOATING
C500 a1 0 0.140495p $ **FLOATING
C501 a_612_n65# 0 44.863f $ **FLOATING
C502 a_924_n35# 0 14.266f $ **FLOATING
C503 a_848_2# 0 31.139002f $ **FLOATING
C504 a_883_n2# 0 3.508f $ **FLOATING
C505 p2 0 0.505775p $ **FLOATING
C506 a_337_67# 0 3.508f $ **FLOATING
C507 a_582_25# 0 18.082f $ **FLOATING
C508 a_879_123# 0 4.916f $ **FLOATING
C509 a_691_36# 0 14.266f $ **FLOATING
C510 a_345_92# 0 14.946f $ **FLOATING
C511 a_302_20# 0 31.139002f $ **FLOATING
C512 a_269_20# 0 14.266f $ **FLOATING
C513 a_324_88# 0 4.916f $ **FLOATING
C514 b0 0 85.82f $ **FLOATING
C515 a0 0 0.144276p $ **FLOATING
C516 s1 0 3.76f $ **FLOATING
C517 c1 0 17.83f $ **FLOATING
C518 a_798_100# 0 14.946f $ **FLOATING
C519 a_615_73# 0 44.863f $ **FLOATING
C520 a_445_140# 0 4.888f $ **FLOATING
C521 a_445_147# 0 20.28f $ **FLOATING
C522 a_907_111# 0 14.266f $ **FLOATING
C523 a_831_148# 0 31.139002f $ **FLOATING
C524 a_866_144# 0 3.508f $ **FLOATING
C525 p1 0 0.380473p $ **FLOATING
C526 pocin 0 28.03f $ **FLOATING
C527 a_271_142# 0 18.082f $ **FLOATING
C528 a_380_153# 0 14.266f $ **FLOATING
C529 a_819_257# 0 4.916f $ **FLOATING
C530 a_496_232# 0 1.316f $ **FLOATING
C531 cin 0 80.576996f $ **FLOATING
C532 p0 0 0.200305p $ **FLOATING
C533 s0 0 3.76f $ **FLOATING
C534 a_738_234# 0 14.946f $ **FLOATING
C535 a_304_190# 0 44.863f $ **FLOATING
C536 a_496_251# 0 1.316f $ **FLOATING
C537 p1p0c0 0 12.783999f $ **FLOATING
C538 a_617_278# 0 4.888f $ **FLOATING
C539 p1g0 0 18.06f $ **FLOATING
C540 a_600_239# 0 21.819f $ **FLOATING
C541 a_847_245# 0 14.266f $ **FLOATING
C542 a_771_282# 0 31.139002f $ **FLOATING
C543 a_806_278# 0 3.508f $ **FLOATING
C544 a_617_318# 0 2.585f $ **FLOATING
C545 g1 0 0.241318p $ **FLOATING
C546 a_453_311# 0 17.907999f $ **FLOATING
C547 a_271_280# 0 18.082f $ **FLOATING
C548 c4 0 4.324f $ **FLOATING
C549 p3p2p1p0c0 0 12.783999f $ **FLOATING
C550 a_380_291# 0 14.266f $ **FLOATING
C551 a_610_377# 0 1.128f $ **FLOATING
C552 g0 0 0.142589p $ **FLOATING
C553 a_304_328# 0 44.863f $ **FLOATING
C554 a_440_393# 0 1.316f $ **FLOATING
C555 a_610_395# 0 1.316f $ **FLOATING
C556 a_883_389# 0 4.888f $ **FLOATING
C557 p3p2p1g0 0 18.624f $ **FLOATING
C558 a_825_350# 0 23.605001f $ **FLOATING
C559 p2g1 0 12.22f $ **FLOATING
C560 a_610_414# 0 1.316f $ **FLOATING
C561 a_440_412# 0 1.316f $ **FLOATING
C562 a_731_417# 0 4.888f $ **FLOATING
C563 p2p1p0c0 0 18.624f $ **FLOATING
C564 a_883_429# 0 2.585f $ **FLOATING
C565 p3p2g1 0 30.286f $ **FLOATING
C566 a_693_378# 0 22.75f $ **FLOATING
C567 a_731_457# 0 2.585f $ **FLOATING
C568 p2p1g0 0 30.286f $ **FLOATING
C569 a_883_464# 0 2.35f $ **FLOATING
C570 p3g2 0 40.25f $ **FLOATING
C571 a_218_418# 0 18.082f $ **FLOATING
C572 a_534_474# 0 18.762999f $ **FLOATING
C573 a_397_472# 0 17.907999f $ **FLOATING
C574 a_327_429# 0 14.266f $ **FLOATING
C575 a_731_492# 0 2.35f $ **FLOATING
C576 g2 0 0.205115p $ **FLOATING
C577 a_884_498# 0 2.115f $ **FLOATING
C578 a_251_466# 0 44.863f $ **FLOATING
C579 a_424_535# 0 1.316f $ **FLOATING
C580 a_594_537# 0 1.316f $ **FLOATING
C581 a_797_547# 0 1.316f $ **FLOATING
C582 a_594_556# 0 1.316f $ **FLOATING
C583 a_424_554# 0 1.316f $ **FLOATING
C584 a_797_566# 0 1.316f $ **FLOATING
C585 a_594_575# 0 1.316f $ **FLOATING
C586 a_797_585# 0 1.316f $ **FLOATING
C587 a_797_604# 0 1.316f $ **FLOATING
C588 a_206_556# 0 18.082f $ **FLOATING
C589 a_315_567# 0 14.266f $ **FLOATING
C590 a_381_614# 0 17.907999f $ **FLOATING
C591 a_239_604# 0 44.863f $ **FLOATING
C592 a_518_635# 0 18.762999f $ **FLOATING
C593 a_688_664# 0 19.618f $ **FLOATING
