* SPICE3 file created from testing.ext - technology: scmos

.option scale=90n

M1000 a_594_537# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1001 a_239_604# p3 g2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_329_n305# a_325_n314# p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 a_218_418# p2 vdd w_205_450# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_825_350# g3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 a_600_239# p1p0c0 a_617_278# w_611_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 s1 p1 c1 w_818_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 c1 a_445_147# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1008 p3p2p1g0 a_518_635# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1009 a_693_378# p2g1 a_731_417# w_725_411# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_564_n251# a2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1011 a_600_239# p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 a_594_n65# a1 b1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 gnd a_269_20# p0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 a_594_556# p2 a_594_537# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 a_445_147# g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1016 a_594_575# p1 a_594_556# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1017 p2g1 a_327_429# vdd w_347_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1018 a_440_412# p1 a_440_393# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_564_n389# a3 vdd w_551_n357# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1020 p1p0c0 a_453_311# vdd w_544_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1021 a3 b3 p3 w_329_n384# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 a_518_635# p3 vdd w_505_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a_731_457# p2p1p0c0 a_731_417# w_725_444# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1024 a_808_n381# p3 vdd w_795_n349# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1025 b2 a2 p2 w_368_n246# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1026 p3p2g1 a_381_614# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 p2p1p0c0 a_534_474# vdd w_658_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1028 a_610_395# p1 a_610_377# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1029 a_329_n171# a_325_n180# p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 a_518_635# g0 a_594_575# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 s2 a_795_n247# a_873_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 vdd a0 a_324_88# w_400_28# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1033 a_594_n65# a_561_n113# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1034 vdd a_302_20# a_269_20# w_291_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 a_325_n180# b2 p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 a_825_350# p3p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1037 a_304_190# a_271_142# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1038 a_847_245# a_771_282# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1039 a_884_498# p3g2 a_883_464# w_878_485# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 a_731_492# p2p1g0 a_731_457# w_725_479# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1041 a_673_n378# a_597_n341# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 a_597_n341# a_564_n389# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1043 a_315_567# a_239_604# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 g0 a_673_36# vdd w_693_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 p3g2 a_315_567# vdd w_335_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 vdd g3 a_884_498# w_879_518# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1047 a_825_350# p3p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 pocin a_380_153# vdd w_400_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 vdd a_269_20# p0 w_258_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 a_218_418# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1051 a_380_153# a_304_190# vdd w_367_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 b1 a1 a_302_n114# w_367_n112# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_825_350# p3p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1054 a_271_280# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1055 p3p2p1g0 a_518_635# vdd w_642_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_239_604# a_206_556# g2 w_226_594# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 a_304_190# a_271_142# cin w_291_180# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 c3 a_693_378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 g3 a_673_n378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 p2p1g0 a_397_472# vdd w_488_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_440_393# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_688_664# p0 vdd w_774_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 s2 p2 c2 w_815_n209# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1064 a_445_147# pocin gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 p2g1 a_327_429# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 a_600_239# p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1067 a_795_n247# p2 vdd w_782_n215# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_564_n251# a2 vdd w_551_n219# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_327_429# a_251_466# vdd w_314_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 a_688_664# cin vdd w_807_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1071 a_693_378# p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_251_466# p2 g1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 s1 c1 a_798_n113# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_798_n113# p1 vdd w_785_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_325_n314# b3 p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 a_738_234# p0 vdd w_725_266# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1077 a_673_36# a_597_73# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1078 a_564_25# a0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1079 p3p2g1 a_381_614# vdd w_472_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1080 a_597_n341# a_564_n389# b3 w_584_n351# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1081 a_206_556# p3 vdd w_193_588# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_424_535# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1083 g2 a_564_n251# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1084 g1 a_670_n102# vdd w_690_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1085 s3 p3 c3 w_828_n343# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_610_377# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1087 s0 a_847_245# vdd w_867_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1088 vdd a2 a_325_n180# w_401_n240# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_670_n102# a_594_n65# vdd w_657_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 c4 a_825_350# vdd w_942_382# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_670_n102# a_594_n65# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_424_554# p2 a_424_535# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 a_453_311# p0 vdd w_473_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1094 a_315_567# a_239_604# vdd w_302_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 p3p2p1p0c0 a_688_664# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_771_282# p0 cin w_758_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1097 s1 c1 p1 w_857_n67# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_271_142# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1099 a_534_474# cin vdd w_620_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_534_474# p0 vdd w_587_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_453_311# cin vdd w_506_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1102 a_271_280# p1 vdd w_258_312# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_561_n113# a1 vdd w_548_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 a_381_614# g1 a_424_554# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_883_429# p3p2p1g0 a_883_389# w_877_416# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_693_378# p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 c1 a_445_147# vdd w_504_133# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_304_328# a_271_280# g0 w_291_318# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 a_825_350# p3g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1110 a_564_n389# a3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 s1 a_798_n113# a_876_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_688_664# p1 vdd w_741_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1113 a_797_604# p0 a_797_585# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 vdd a_269_n114# p1 w_258_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1115 p1g0 a_380_291# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_324_n46# b1 a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 a_327_429# a_251_466# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1118 a_693_378# p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 a_380_291# a_304_328# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1120 c2 a_600_239# vdd w_676_271# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 b3 a3 p3 w_368_n380# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1122 a1 b1 a_302_n114# w_328_n116# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 a_328_n37# a_324_n46# a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1124 a_328_97# a_324_88# a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 vdd a3 a_325_n314# w_401_n374# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1126 a_597_n341# a3 b3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 p1p0c0 a_453_311# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1128 a_324_88# b0 a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1129 a_688_664# cin a_797_604# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 vdd g2 a_731_492# w_726_513# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1131 a_883_464# p3p2g1 a_883_429# w_877_451# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_693_378# g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_304_328# p1 g0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1134 g2 a_564_n251# b2 w_584_n213# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1135 a_597_73# a_564_25# b0 w_584_63# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1136 a_597_73# a0 b0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1137 a_771_282# a_738_234# a_816_233# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1138 a_518_635# p1 vdd w_571_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_397_472# g0 vdd w_450_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_797_547# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_496_251# p0 a_496_232# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 a_847_245# a_771_282# vdd w_834_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_597_73# a_564_25# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1147 a_239_604# a_206_556# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1148 a_797_566# p2 a_797_547# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1149 a_453_311# cin a_496_251# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1150 a_453_311# p1 vdd w_440_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 gnd a3 a_325_n314# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1152 a_534_474# p1 vdd w_554_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_304_328# a_271_280# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1154 a_445_147# g0 a_445_140# w_439_134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 a_797_585# p1 a_797_566# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 gnd a_302_n114# a_269_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_795_n247# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1158 gnd a_269_n114# p1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1159 g0 a_673_36# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1160 a_381_614# g1 vdd w_434_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 s2 c2 a_795_n247# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_561_n113# a1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1163 pocin a_380_153# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_380_153# a_304_190# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1165 a_688_664# p3 vdd w_675_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1166 s3 a_808_n381# a_886_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1167 a_673_n378# a_597_n341# vdd w_660_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 g2 a2 b2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 p1g0 a_380_291# vdd w_400_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1170 c2 a_600_239# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 g1 a_670_n102# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1172 a0 b0 a_302_20# w_328_18# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 a_380_291# a_304_328# vdd w_367_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_688_664# p2 vdd w_708_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1175 p2p1g0 a_397_472# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1176 gnd a2 a_325_n180# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 vdd pocin a_445_140# w_439_167# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1178 c3 a_693_378# vdd w_790_410# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_304_190# p0 cin Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1180 s3 c3 a_808_n381# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1181 a_251_466# a_218_418# g1 w_238_456# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1182 s3 c3 p3 w_867_n335# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 vdd a1 a_324_n46# w_400_n106# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1184 a_673_36# a_597_73# vdd w_660_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1185 a_397_472# g0 a_440_412# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 a_808_n381# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1187 a_798_n113# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_564_25# a0 vdd w_551_57# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 g3 a_673_n378# vdd w_693_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# p2 vdd w_384_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 vdd a_302_n114# a_269_n114# w_291_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1192 a_617_318# p1g0 a_617_278# w_611_305# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1193 a_771_282# cin p0 w_797_280# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 a_738_234# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1195 a_594_n65# a_561_n113# b1 w_581_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_518_635# p2 vdd w_538_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 b0 a0 a_302_20# w_367_22# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_496_232# p1 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1199 a_397_472# p1 vdd w_417_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_206_556# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1201 p3p2p1p0c0 a_688_664# vdd w_845_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 a_610_414# p0 a_610_395# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_534_474# p2 vdd w_521_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_271_142# p0 vdd w_258_174# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1205 s0 a_847_245# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 vdd g1 a_617_318# w_611_340# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 c4 a_825_350# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1208 gnd a1 a_324_n46# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1209 gnd a0 a_324_88# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 gnd a_302_20# a_269_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1211 a_381_614# p2 vdd w_401_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1212 a2 b2 p2 w_329_n250# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 a_251_466# a_218_418# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 a_534_474# cin a_610_414# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1215 a_771_282# cin a_738_234# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 a_381_614# p3 vdd w_368_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1217 p3g2 a_315_567# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1218 a_600_239# g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1219 s2 c2 p2 w_854_n201# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 w_725_411# a_693_378# 0.013329f
C1 p3g2 w_878_485# 0.036563f
C2 p3p2p1g0 w_879_518# 0.011197f
C3 p2p1p0c0 p2p1g0 0.049073f
C4 p3p2g1 g0 0.011924f
C5 g1 p1p0c0 0.002848f
C6 g2 p3 0.016679f
C7 g3 p1 0.028063f
C8 a0 p0 0.007627f
C9 a_771_282# gnd 0.190422f
C10 p0 c2 0.020959f
C11 w_867_277# s0 0.013216f
C12 g0 p2g1 0.002352f
C13 a_797_566# p2 0.013746f
C14 a_424_554# p3 0.025115f
C15 a_381_614# w_401_604# 0.027639f
C16 w_258_312# vdd 0.0086f
C17 a_731_492# vdd 0.41238f
C18 g3 gnd 0.214319f
C19 p3 p0 0.002576f
C20 w_693_68# vdd 0.008451f
C21 a_825_350# w_942_382# 0.027289f
C22 a_883_389# w_877_383# 0.017071f
C23 p2 p1 2.60374f
C24 a_271_280# vdd 0.439891f
C25 w_258_174# p0 0.028034f
C26 b1 a_328_n37# 0.001802f
C27 a_302_20# vdd 0.019283f
C28 w_725_266# c2 0.003448f
C29 p2g1 w_384_462# 1.09e-20
C30 c4 a_825_350# 0.060798f
C31 a_397_472# w_488_462# 0.027163f
C32 b0 gnd 0.035498f
C33 a_324_n46# a_302_n114# 0.286223f
C34 vdd s0 0.439883f
C35 a_302_20# w_291_17# 0.027261f
C36 c3 s0 0.003003f
C37 w_439_167# pocin 0.036563f
C38 a_327_429# p2g1 0.060798f
C39 g2 a_564_n251# 0.003752f
C40 a_594_n65# a_670_n102# 0.060798f
C41 cin vdd 0.044543f
C42 p2 gnd 1.792362f
C43 a_251_466# w_238_456# 0.019526f
C44 c3 cin 5.08e-19
C45 c1 w_504_133# 0.013242f
C46 c2 a_873_n248# 0.001866f
C47 w_367_185# a_304_190# 0.026907f
C48 w_544_301# g0 0.00229f
C49 w_611_340# g1 0.039692f
C50 a_731_492# p2p1g0 3.63e-19
C51 g1 vdd 0.773639f
C52 p3 w_329_n384# 0.007992f
C53 p2 w_854_n201# 0.007896f
C54 p3 a_325_n314# 0.286223f
C55 w_758_272# vdd 6.13e-19
C56 p3p2p1p0c0 a_688_664# 0.060798f
C57 p3p2p1g0 a_518_635# 0.060798f
C58 a_797_604# cin 0.013759f
C59 a_594_575# p1 0.031835f
C60 a_797_585# p0 0.013746f
C61 p2 s2 0.413834f
C62 a_808_n381# a_886_n382# 0.14502f
C63 a_304_328# vdd 0.017291f
C64 w_329_n250# p2 0.011491f
C65 w_741_654# a_688_664# 0.027639f
C66 w_205_450# p2 0.028034f
C67 w_857_n67# p1 0.007896f
C68 w_328_n116# b1 0.027716f
C69 w_367_n112# a1 0.028748f
C70 a_884_498# w_878_485# 0.01128f
C71 w_258_n117# a_269_n114# 0.026907f
C72 a_424_554# a_381_614# 0.41238f
C73 a_251_466# a_218_418# 0.003752f
C74 a_798_n113# c2 0.003242f
C75 cin p2p1g0 3.55e-20
C76 p3g2 p3 0.026608f
C77 g2 w_193_588# 0.009535f
C78 w_551_n357# a3 0.02808f
C79 w_584_n351# a_597_n341# 0.019526f
C80 a_564_n389# a3 0.060856f
C81 gnd a_795_n247# 0.206673f
C82 vdd a_597_n341# 0.011738f
C83 a_445_140# pocin 0.185571f
C84 w_401_n240# vdd 0.008451f
C85 cin w_620_464# 0.026794f
C86 p1 a_670_n102# 0.002494f
C87 p0 g0 0.011127f
C88 p2 a_534_474# 0.002444f
C89 p1 a_397_472# 0.017711f
C90 a_693_378# gnd 1.08291f
C91 w_815_n209# s2 0.015055f
C92 a_315_567# gnd 0.248155f
C93 p3p2g1 vdd 0.439963f
C94 p1 w_571_625# 0.026996f
C95 p1p0c0 w_544_301# 0.013229f
C96 vdd a2 0.195509f
C97 p1p0c0 a_600_239# 0.211061f
C98 p3g2 a_825_350# 0.001345f
C99 a_795_n247# s2 0.286223f
C100 w_581_n75# vdd 2.04e-19
C101 w_675_654# vdd 0.008451f
C102 a_771_282# a_816_233# 0.20619f
C103 p1 w_417_462# 0.026996f
C104 pocin a_445_147# 1.39e-20
C105 a_670_n102# gnd 0.248155f
C106 w_790_410# vdd 0.008451f
C107 c3 s1 0.003481f
C108 p2g1 vdd 0.439883f
C109 a_397_472# gnd 0.042086f
C110 c3 w_790_410# 0.013216f
C111 p3g2 a_797_585# 0.054573f
C112 g3 a_771_282# 2.33e-19
C113 p3p2g1 a_797_604# 0.003102f
C114 p3 w_368_604# 0.026794f
C115 p3p2p1g0 p3p2p1p0c0 0.003212f
C116 a_440_393# g0 7.76e-19
C117 c3 a_876_n114# 6.44e-19
C118 b2 a_325_n180# 0.02927f
C119 g1 w_347_461# 0.01132f
C120 a_673_36# w_693_68# 0.026907f
C121 vdd w_521_464# 0.008451f
C122 b1 vdd 0.015576f
C123 p3p2p1g0 w_877_416# 0.03763f
C124 p3p2p1p0c0 w_877_451# 0.018013f
C125 a_381_614# p3g2 0.011947f
C126 p3p2p1g0 a_883_464# 0.016011f
C127 p1 w_440_301# 0.026794f
C128 w_439_167# g0 4.29e-19
C129 g2 a_239_604# 0.75303f
C130 vdd w_401_604# 0.008451f
C131 a_453_311# cin 0.069062f
C132 a_597_73# w_660_68# 0.026907f
C133 a_324_88# w_400_28# 0.013216f
C134 a_564_25# p0 0.003966f
C135 cin a_380_153# 0.003392f
C136 a0 a_324_88# 0.060798f
C137 p0 a_271_142# 0.060798f
C138 w_877_451# a_883_464# 0.01128f
C139 p3p2g1 w_879_518# 4.09e-19
C140 a_594_556# a_594_537# 0.41238f
C141 a_424_554# a_424_535# 0.41238f
C142 p2g1 p2p1g0 0.005273f
C143 p3g2 g0 7.61e-19
C144 g3 p2 0.022389f
C145 w_544_301# vdd 0.008451f
C146 a_304_328# w_367_323# 0.026907f
C147 a_600_239# vdd 0.001532f
C148 a_597_73# p0 0.007562f
C149 p1 c2 0.003604f
C150 gnd pocin 0.372676f
C151 g3 w_693_n346# 0.013222f
C152 w_942_382# vdd 0.008451f
C153 c1 g1 0.008592f
C154 a_315_567# w_335_599# 0.026907f
C155 a_381_614# w_368_604# 0.017642f
C156 g2 vdd 0.029171f
C157 a_251_466# gnd 0.701773f
C158 p3 p1 0.040972f
C159 a_825_350# w_877_383# 0.013329f
C160 w_660_68# vdd 0.008507f
C161 c4 vdd 0.439883f
C162 b1 a_302_n114# 0.685112f
C163 a_269_20# vdd 0.441416f
C164 p2g1 w_347_461# 0.013223f
C165 w_676_271# c2 0.016933f
C166 a_397_472# w_450_462# 0.027639f
C167 a0 gnd 1.211792f
C168 vdd a_738_234# 0.439891f
C169 gnd c2 0.219293f
C170 b0 w_367_22# 0.01395f
C171 a_269_20# w_291_17# 0.013216f
C172 w_400_185# pocin 0.013216f
C173 a_445_140# g0 0.016231f
C174 g2 w_584_n213# 0.019526f
C175 w_611_340# p0 4.94e-20
C176 p0 vdd 0.73653f
C177 p3 gnd 1.577599f
C178 w_854_n201# c2 0.027735f
C179 a_610_414# cin 0.013746f
C180 c3 p0 1.47e-20
C181 c2 s2 0.686118f
C182 w_291_180# a_304_190# 0.019526f
C183 a_797_566# a_797_585# 0.41238f
C184 p2 w_815_n209# 0.028748f
C185 p3p2g1 a_518_635# 0.041586f
C186 p3 b3 0.685112f
C187 a_797_604# p0 0.013746f
C188 p3p2p1g0 a_688_664# 0.00431f
C189 a_797_585# p1 0.013746f
C190 w_725_266# vdd 0.0086f
C191 p2 a_795_n247# 0.060798f
C192 g0 a_445_147# 0.216537f
C193 a_808_n381# gnd 0.206673f
C194 c3 a_886_n382# 0.002154f
C195 a_825_350# gnd 1.35993f
C196 w_818_n75# p1 0.028748f
C197 w_774_654# p0 0.026996f
C198 w_708_654# a_688_664# 0.027639f
C199 a_731_492# w_726_513# 0.009864f
C200 w_328_n116# a1 0.007896f
C201 c1 s1 0.686034f
C202 a_380_291# g0 0.008577f
C203 a_206_556# p3 0.069923f
C204 p0 p2p1g0 0.001001f
C205 c1 a_876_n114# 0.001856f
C206 g1 w_690_n70# 0.01323f
C207 a_325_n314# vdd 0.439883f
C208 w_401_n374# a3 0.028034f
C209 a_564_n389# a_597_n341# 0.003752f
C210 gnd a_564_n251# 0.20619f
C211 w_439_167# vdd 0.010186f
C212 c3 a_873_n248# 4.29e-20
C213 w_238_456# vdd 6.13e-19
C214 p1 a_328_n37# 6.43e-21
C215 cin w_726_513# 0.002754f
C216 p2 a_397_472# 0.002835f
C217 p1 g0 0.057312f
C218 a_453_311# w_544_301# 0.027163f
C219 p3g2 vdd 0.440124f
C220 a_381_614# gnd 0.042086f
C221 p1g0 a_617_278# 0.004158f
C222 w_548_n81# vdd 0.0086f
C223 w_642_625# vdd 0.008451f
C224 w_401_n240# a_325_n180# 0.013216f
C225 a_798_n113# vdd 0.439883f
C226 c3 a_798_n113# 0.001329f
C227 a_380_291# w_400_323# 0.026907f
C228 a_218_418# vdd 0.439891f
C229 g0 gnd 0.208112f
C230 a_271_280# w_291_318# 0.026794f
C231 p3p2g1 p3p2p1p0c0 0.001238f
C232 p3p2p1p0c0 a_883_429# 0.005194f
C233 a_610_414# p2g1 0.019171f
C234 g1 w_314_461# 0.01132f
C235 a2 a_325_n180# 0.060798f
C236 a_673_36# w_660_68# 0.013216f
C237 a_564_25# w_584_63# 0.026794f
C238 a_302_20# a_328_97# 0.20619f
C239 a_771_282# c2 0.020436f
C240 vdd w_488_462# 0.008451f
C241 c2 a_816_233# 3.8e-19
C242 a_304_190# a_271_142# 0.003752f
C243 a1 vdd 0.229007f
C244 a_883_429# w_877_416# 0.009864f
C245 p3p2p1g0 w_877_451# 0.012016f
C246 a_327_429# gnd 0.248155f
C247 p3p2g1 a_883_464# 3.63e-19
C248 a_883_429# a_883_464# 0.41238f
C249 w_785_n81# a_798_n113# 0.013216f
C250 a_445_140# vdd 0.41238f
C251 a_597_73# w_584_63# 0.019526f
C252 b0 w_400_28# 0.015139f
C253 p1g0 cin 0.012177f
C254 a_453_311# p0 0.005763f
C255 a0 w_551_57# 0.028093f
C256 vdd w_368_604# 0.008451f
C257 w_867_277# a_847_245# 0.026907f
C258 g3 c2 0.005387f
C259 a0 b0 0.539271f
C260 a_673_36# p0 0.003088f
C261 cin a_496_232# 0.024151f
C262 a_594_n65# vdd 0.013824f
C263 w_725_444# a_731_457# 0.009864f
C264 g1 p1g0 0.038781f
C265 a_251_466# p2 0.001371f
C266 a_797_547# cin 2.48e-20
C267 w_506_301# vdd 0.008451f
C268 p3p2g1 w_472_604# 0.013216f
C269 w_604_625# g0 0.026794f
C270 a_206_556# w_193_588# 0.013216f
C271 a_304_328# w_291_318# 0.019526f
C272 cin a_688_664# 0.059029f
C273 a_847_245# vdd 0.441416f
C274 c1 p0 0.015446f
C275 p1p0c0 gnd 0.207724f
C276 a_847_245# c3 0.006337f
C277 p2 c2 0.026943f
C278 a_564_25# gnd 0.20619f
C279 p2p1g0 w_488_462# 0.013216f
C280 gnd a_271_142# 0.20619f
C281 vdd a_445_147# 0.001532f
C282 w_658_464# p2p1p0c0 0.013216f
C283 a_315_567# w_302_599# 0.013216f
C284 a_424_535# gnd 0.41238f
C285 a_884_498# vdd 0.41238f
C286 g3 a_825_350# 0.002823f
C287 p3 p2 0.395341f
C288 w_584_63# vdd 2.04e-19
C289 a_380_291# vdd 0.441416f
C290 w_797_280# cin 0.027729f
C291 a_239_604# gnd 0.248155f
C292 a_324_88# vdd 0.439891f
C293 g0 w_450_462# 0.026794f
C294 a_397_472# w_417_462# 0.027639f
C295 a_597_73# gnd 0.248155f
C296 a1 a_302_n114# 0.413834f
C297 vdd a_304_190# 0.017997f
C298 a_269_20# w_258_17# 0.026907f
C299 b0 w_328_18# 0.027757f
C300 a0 w_367_22# 0.028748f
C301 p3 s3 0.413834f
C302 p1 vdd 0.832418f
C303 w_815_n209# c2 0.01623f
C304 w_258_17# p0 0.013216f
C305 a_610_414# p0 0.019134f
C306 c2 a_795_n247# 0.017003f
C307 p2 w_782_n215# 0.028034f
C308 p3p2p1g0 cin 0.02473f
C309 a_206_556# a_239_604# 0.003752f
C310 a_594_575# p3 2.95e-20
C311 p3g2 a_518_635# 8.1e-19
C312 w_611_340# gnd 1.17e-19
C313 w_676_271# vdd 0.008451f
C314 p2 a_564_n251# 0.002692f
C315 vdd gnd 2.215753f
C316 a_808_n381# s3 0.286223f
C317 c3 gnd 0.223819f
C318 w_642_625# a_518_635# 0.027163f
C319 a_825_350# a_883_389# 0.453641f
C320 w_785_n81# p1 0.028309f
C321 w_675_654# a_688_664# 0.017642f
C322 a_884_498# w_879_518# 0.009864f
C323 g2 w_726_513# 0.036563f
C324 c1 a_798_n113# 0.016996f
C325 g3 g0 0.00202f
C326 g1 b2 7.83e-19
C327 a_315_567# p3 0.001362f
C328 a_381_614# p2 0.005763f
C329 cin p2p1p0c0 0.007704f
C330 p1 p2p1g0 0.008846f
C331 b3 w_584_n351# 0.008451f
C332 b3 vdd 0.013251f
C333 w_368_n380# a3 0.028748f
C334 c3 w_854_n201# 5.29e-20
C335 a_673_n378# a_597_n341# 0.060798f
C336 w_400_185# vdd 0.008451f
C337 a_597_n341# a3 0.001371f
C338 c3 s2 0.015855f
C339 w_205_450# vdd 0.0086f
C340 p0 w_587_464# 0.026996f
C341 p1 a_302_n114# 0.007287f
C342 p2 g0 0.033881f
C343 a_453_311# w_506_301# 0.027639f
C344 p1g0 w_544_301# 0.004305f
C345 p2p1g0 gnd 0.207724f
C346 w_782_n215# a_795_n247# 0.013216f
C347 a_206_556# vdd 0.439891f
C348 p2 w_538_625# 0.026794f
C349 p1g0 a_600_239# 0.040556f
C350 w_604_625# vdd 0.008451f
C351 p2 w_384_462# 0.026794f
C352 w_551_n219# a2 0.028079f
C353 w_401_n240# b2 0.015139f
C354 a_302_n114# gnd 0.190422f
C355 a_561_n113# vdd 0.439891f
C356 g1 w_434_604# 0.026794f
C357 a_534_474# vdd 1.76176f
C358 a_271_280# w_258_312# 0.013216f
C359 a_380_291# w_367_323# 0.013216f
C360 p3g2 p3p2p1p0c0 0.001239f
C361 p3p2g1 p3p2p1g0 0.0533f
C362 a_731_417# p2p1p0c0 0.004158f
C363 p3p2p1g0 a_883_429# 0.00801f
C364 a_564_25# w_551_57# 0.013216f
C365 a2 b2 0.531092f
C366 b0 a_564_25# 0.00288f
C367 c1 a_445_147# 0.060798f
C368 vdd w_450_462# 0.008451f
C369 a_304_190# a_380_153# 0.060798f
C370 p3p2g1 w_877_451# 0.037044f
C371 a_883_429# w_877_451# 0.009864f
C372 a_594_575# g0 0.013746f
C373 p1g0 p0 7.17e-19
C374 a0 w_400_28# 0.028034f
C375 vdd w_335_599# 0.008451f
C376 a_453_311# p1 0.002444f
C377 w_834_277# a_847_245# 0.013216f
C378 a_328_97# p0 3.98e-19
C379 a_597_73# b0 0.756776f
C380 p0 a_496_232# 0.013746f
C381 p2g1 p2p1p0c0 0.008706f
C382 a_424_535# p2 0.023137f
C383 w_473_301# vdd 0.008451f
C384 w_611_272# p1p0c0 0.057514f
C385 w_611_305# a_617_318# 0.009864f
C386 w_400_n106# vdd 0.0086f
C387 c1 p1 0.024407f
C388 p1 a_518_635# 0.005763f
C389 p0 a_688_664# 0.005763f
C390 a_453_311# gnd 0.042086f
C391 a_771_282# vdd 0.019283f
C392 a_771_282# c3 0.007917f
C393 a_271_280# a_304_328# 0.003752f
C394 a_534_474# w_620_464# 0.027639f
C395 a_673_36# gnd 0.248155f
C396 gnd a_380_153# 0.248155f
C397 g0 a_397_472# 0.059421f
C398 g1 cin 0.016729f
C399 a_594_537# gnd 0.41238f
C400 g3 vdd 0.446831f
C401 w_797_280# p0 0.007968f
C402 w_758_272# cin 0.013523f
C403 w_551_57# vdd 0.0086f
C404 g2 a3 0.009821f
C405 g3 c3 0.073145f
C406 a_518_635# gnd 0.042086f
C407 a_610_377# p0 6.84e-20
C408 b1 a_324_n46# 0.02927f
C409 a_397_472# w_384_462# 0.017642f
C410 c1 gnd 0.206382f
C411 b0 vdd 0.015588f
C412 a0 w_328_18# 0.007896f
C413 w_400_185# a_380_153# 0.026907f
C414 g2 w_226_594# 0.018971f
C415 p3p2p1p0c0 w_877_383# 0.053825f
C416 a_884_498# p3p2p1p0c0 0.005507f
C417 g2 b2 0.764942f
C418 p3 a_808_n381# 0.060798f
C419 w_867_n335# s3 0.007992f
C420 p2 vdd 0.639134f
C421 w_818_n75# c2 0.019549f
C422 a_884_498# a_883_464# 0.41238f
C423 a_797_547# p3g2 0.001272f
C424 g2 p2p1p0c0 0.063553f
C425 p3p2g1 cin 0.004802f
C426 p3p2p1g0 p0 0.013798f
C427 a_315_567# a_239_604# 0.060798f
C428 vdd w_693_n346# 0.008451f
C429 a_564_n389# gnd 0.20619f
C430 p2 a_329_n171# 0.20619f
C431 c3 s3 0.692464f
C432 a_440_412# a_440_393# 0.41238f
C433 a_610_414# a_610_395# 0.41238f
C434 w_604_625# a_518_635# 0.027639f
C435 w_367_22# vdd 6.13e-19
C436 w_690_n70# p1 0.002922f
C437 w_741_654# p1 0.026794f
C438 g3 w_879_518# 0.036563f
C439 g1 a2 0.011016f
C440 p0 p2p1p0c0 0.002479f
C441 cin p2g1 0.013147f
C442 p2 p2p1g0 7.61e-20
C443 a_381_614# p3 0.003255f
C444 a_325_n314# w_401_n374# 0.013216f
C445 b3 a_564_n389# 0.00288f
C446 w_329_n384# a3 0.007896f
C447 p3p2p1p0c0 gnd 0.207724f
C448 vdd a_795_n247# 0.439891f
C449 gnd a_325_n180# 0.206673f
C450 a_325_n314# a3 0.060798f
C451 w_367_185# vdd 0.008465f
C452 c3 a_795_n247# 4.01e-19
C453 a_600_239# a_617_278# 0.453641f
C454 w_845_654# vdd 0.008451f
C455 a_251_466# a_327_429# 0.060798f
C456 p1 a_269_n114# 0.06333f
C457 g1 p2g1 0.007851f
C458 p1g0 w_506_301# 0.004305f
C459 a_693_378# vdd 0.001532f
C460 a_453_311# w_473_301# 0.027639f
C461 a_315_567# vdd 0.441416f
C462 a_239_604# w_302_599# 0.026907f
C463 w_193_588# p3 0.028034f
C464 c3 a_693_378# 0.060798f
C465 g1 b1 0.281479f
C466 w_368_n246# b2 0.01395f
C467 w_401_n240# a2 0.028034f
C468 a_670_n102# vdd 0.441416f
C469 a_269_n114# gnd 0.248155f
C470 a_397_472# vdd 1.32165f
C471 p3g2 p3p2p1g0 0.001431f
C472 a_610_414# a_534_474# 0.41238f
C473 a_731_417# p2g1 0.019622f
C474 a_380_291# p1g0 0.060798f
C475 vdd w_571_625# 0.008451f
C476 a_600_239# cin 8.95e-19
C477 a_453_311# a_496_251# 0.41238f
C478 p3p2p1g0 w_642_625# 0.013284f
C479 a_324_88# a_328_97# 0.14502f
C480 a_269_20# a_302_20# 0.060798f
C481 a0 a_564_25# 0.060867f
C482 vdd w_417_462# 0.008451f
C483 p2p1g0 a_693_378# 0.001345f
C484 g1 a_600_239# 1.39e-20
C485 g2 cin 0.003885f
C486 w_258_n117# p1 0.013216f
C487 w_693_68# p0 0.001671f
C488 c1 g3 0.003696f
C489 vdd w_302_599# 0.008507f
C490 p1g0 p1 7.17e-19
C491 w_834_277# a_771_282# 0.027261f
C492 a_302_20# p0 0.003749f
C493 a_597_73# a0 0.001371f
C494 cin a_738_234# 0.024367f
C495 w_258_174# a_271_142# 0.013216f
C496 p1 a_496_232# 0.013746f
C497 s1 a_876_n114# 0.20619f
C498 w_725_479# a_731_457# 0.009864f
C499 w_725_411# p2p1p0c0 0.001174f
C500 a_797_566# a_797_547# 0.41238f
C501 g2 g1 1.63579f
C502 a_397_472# p2p1g0 0.060798f
C503 a_594_537# p2 0.020283f
C504 a_424_535# p3 0.013746f
C505 w_581_n75# b1 0.009938f
C506 w_834_277# g3 0.016049f
C507 w_440_301# vdd 0.008451f
C508 w_611_340# a_617_318# 0.009864f
C509 p3 a_239_604# 0.002112f
C510 p0 cin 0.261159f
C511 w_611_305# p1p0c0 1.04e-20
C512 p1 a_688_664# 0.004034f
C513 p2 a_518_635# 0.004034f
C514 w_367_n112# vdd 6.13e-19
C515 a_617_318# vdd 0.41238f
C516 p1g0 gnd 0.207724f
C517 a_534_474# w_587_464# 0.027639f
C518 gnd a_496_232# 0.41238f
C519 vdd pocin 0.439883f
C520 w_504_133# a_445_147# 0.027289f
C521 a_424_554# g1 0.013746f
C522 w_657_n70# a_594_n65# 0.026907f
C523 g1 p0 0.031532f
C524 a_251_466# vdd 0.017997f
C525 w_867_n335# p3 0.007896f
C526 a_797_547# gnd 0.41238f
C527 w_758_272# p0 0.028748f
C528 g2 a_597_n341# 0.013288f
C529 w_400_28# vdd 0.0086f
C530 a1 a_324_n46# 0.060798f
C531 a_688_664# gnd 0.042086f
C532 a_610_377# p1 0.013746f
C533 a0 vdd 0.234154f
C534 vdd c2 0.442422f
C535 c3 c2 0.026004f
C536 w_291_180# a_271_142# 0.026794f
C537 w_367_185# a_380_153# 0.013216f
C538 p3p2p1g0 w_877_383# 0.001142f
C539 a_884_498# p3p2p1g0 0.016011f
C540 g3 p3p2p1p0c0 0.001229f
C541 g2 a2 0.012963f
C542 a_594_575# a_518_635# 0.41238f
C543 p3 vdd 0.976896f
C544 w_828_n343# s3 0.015055f
C545 a_440_412# p1 0.013746f
C546 w_258_174# vdd 0.0086f
C547 c3 p3 0.028649f
C548 a_610_377# gnd 0.41238f
C549 a_610_395# a_610_377# 0.41238f
C550 c1 w_857_n67# 0.027735f
C551 w_367_n112# a_302_n114# 0.015055f
C552 g2 p2g1 0.002942f
C553 w_400_323# g0 0.011443f
C554 p1p0c0 g0 0.010775f
C555 p3p2p1g0 p1 0.010267f
C556 p3p2g1 p0 0.0124f
C557 p3g2 cin 0.004802f
C558 vdd w_660_n346# 0.008507f
C559 p2 a_325_n180# 0.288532f
C560 vdd a_808_n381# 0.439891f
C561 a_673_n378# gnd 0.248155f
C562 g1 w_238_456# 0.021496f
C563 c3 a_808_n381# 0.017003f
C564 w_328_18# vdd 0.001288f
C565 a_825_350# vdd 0.001532f
C566 gnd a3 0.414526f
C567 w_657_n70# p1 0.002922f
C568 c3 a_825_350# 2.29e-19
C569 g1 p3g2 0.023512f
C570 p0 p2g1 0.00813f
C571 vdd w_782_n215# 0.008518f
C572 b3 w_401_n374# 0.015139f
C573 a_325_n314# a_329_n305# 0.14502f
C574 p3p2p1g0 gnd 0.223584f
C575 a_518_635# w_571_625# 0.027639f
C576 b3 a3 0.535308f
C577 w_291_180# vdd 6.13e-19
C578 p3p2p1p0c0 a_883_389# 0.016619f
C579 vdd a_564_n251# 0.439891f
C580 gnd b2 0.037864f
C581 w_807_654# vdd 0.008451f
C582 p1 w_554_464# 0.041309f
C583 p1 a_324_n46# 0.008083f
C584 g1 a_218_418# 0.012164f
C585 a_381_614# vdd 1.32165f
C586 w_584_n213# a_564_n251# 0.026794f
C587 p1g0 w_473_301# 0.004305f
C588 p2p1p0c0 gnd 0.207724f
C589 a_883_389# w_877_416# 0.008113f
C590 a_453_311# w_440_301# 0.017642f
C591 p3 w_505_625# 0.026794f
C592 a_797_604# a_797_585# 0.41238f
C593 a_847_245# s0 0.060798f
C594 p3p2p1p0c0 w_845_654# 0.013216f
C595 g1 a1 0.115698f
C596 w_368_n246# a2 0.028748f
C597 w_329_n250# b2 0.027716f
C598 a_380_153# pocin 0.060798f
C599 a_324_n46# gnd 0.206673f
C600 a_206_556# w_226_594# 0.026794f
C601 a_731_417# w_725_411# 0.017071f
C602 c4 w_942_382# 0.013216f
C603 g0 vdd 0.562964f
C604 cin w_506_301# 0.026794f
C605 p3g2 p3p2g1 0.633236f
C606 vdd w_538_625# 0.008451f
C607 w_193_588# vdd 0.0086f
C608 a_597_73# a_564_25# 0.003752f
C609 b0 a_328_97# 0.001802f
C610 a_324_88# a_302_20# 0.286223f
C611 a_496_251# a_496_232# 0.41238f
C612 vdd w_384_462# 0.008451f
C613 p3p2p1p0c0 w_878_485# 0.018136f
C614 a_327_429# vdd 0.441416f
C615 p1 w_258_312# 0.028034f
C616 g2 p0 0.003358f
C617 w_690_n70# a_670_n102# 0.026907f
C618 w_660_68# p0 0.004686f
C619 a_271_280# p1 0.060798f
C620 a_445_140# w_439_134# 0.017071f
C621 w_797_280# a_771_282# 0.007992f
C622 a_269_20# p0 0.06476f
C623 cin a_304_190# 0.747651f
C624 p0 a_738_234# 0.060798f
C625 a_798_n113# s1 0.286223f
C626 c1 c2 0.013027f
C627 w_725_411# p2g1 0.049155f
C628 w_878_485# a_883_464# 0.009864f
C629 w_725_479# p2p1g0 0.036563f
C630 a_798_n113# a_876_n114# 0.14502f
C631 w_725_444# p2p1p0c0 0.036782f
C632 a_534_474# p2p1p0c0 0.060798f
C633 a_797_566# cin 2.14e-20
C634 a_797_547# p2 0.013746f
C635 a_594_537# p3 0.013776f
C636 a_594_556# p1 0.018694f
C637 w_400_323# vdd 0.008451f
C638 p2 a_688_664# 0.004034f
C639 w_611_272# p1g0 0.001158f
C640 p3 a_518_635# 0.002444f
C641 p1 cin 0.034484f
C642 a_271_280# gnd 0.20619f
C643 p1p0c0 vdd 0.439883f
C644 w_328_n116# vdd 0.001288f
C645 a_380_291# a_304_328# 0.060798f
C646 a_302_n114# a_328_n37# 0.20619f
C647 w_834_277# c2 8.35e-21
C648 w_725_266# a_738_234# 0.013216f
C649 a_302_20# gnd 0.190422f
C650 a_534_474# w_554_464# 0.027639f
C651 a_564_25# vdd 0.439891f
C652 vdd a_271_142# 0.439891f
C653 gnd s0 0.20619f
C654 w_439_134# a_445_147# 0.013329f
C655 w_658_464# a_534_474# 0.027163f
C656 w_581_n75# a_594_n65# 0.019526f
C657 g1 p1 0.015873f
C658 g3 a_673_n378# 0.060798f
C659 w_828_n343# p3 0.028748f
C660 w_725_266# p0 0.028034f
C661 a1 b1 0.614689f
C662 a_239_604# vdd 0.017997f
C663 cin gnd 0.058266f
C664 a_597_73# vdd 0.013824f
C665 a_610_377# p2 0.013746f
C666 a_304_328# p1 0.04464f
C667 w_676_271# g1 0.002127f
C668 g3 p3p2p1g0 0.001198f
C669 g1 gnd 0.373308f
C670 a_327_429# w_347_461# 0.026907f
C671 a_594_n65# b1 0.7623f
C672 w_867_277# vdd 0.008451f
C673 a_440_412# p2 0.011867f
C674 c3 w_867_n335# 0.027759f
C675 w_867_277# c3 3.18e-20
C676 w_400_185# cin 0.00869f
C677 a_304_328# gnd 0.588369f
C678 w_845_654# a_688_664# 0.027163f
C679 c1 w_818_n75# 0.015306f
C680 w_400_n106# a_324_n46# 0.013216f
C681 w_328_n116# a_302_n114# 0.007992f
C682 w_367_323# g0 0.011382f
C683 p3g2 p0 0.002921f
C684 p3p2p1g0 p2 0.010267f
C685 a_673_36# g0 0.060812f
C686 p3p2g1 p1 0.017215f
C687 p2 b2 0.6987f
C688 w_611_340# vdd 0.013119f
C689 a_673_n378# w_693_n346# 0.026907f
C690 g1 w_205_450# 0.013044f
C691 c3 vdd 0.446487f
C692 w_291_17# vdd 0.008507f
C693 gnd a_597_n341# 0.701773f
C694 w_708_654# p2 0.026794f
C695 w_581_n75# p1 0.002922f
C696 p1 s1 0.413834f
C697 a_518_635# g0 0.059018f
C698 p1 p2g1 0.03968f
C699 cin a_534_474# 0.061353f
C700 c1 g0 0.031415f
C701 b3 w_368_n380# 0.01395f
C702 b3 a_329_n305# 0.001802f
C703 p3p2g1 gnd 0.224641f
C704 a_518_635# w_538_625# 0.027639f
C705 p3p2p1p0c0 a_825_350# 0.217915f
C706 b3 a_597_n341# 0.756931f
C707 gnd a2 1.559369f
C708 p3p2p1g0 a_883_389# 0.004158f
C709 a_251_466# w_314_461# 0.026907f
C710 w_785_n81# vdd 0.008451f
C711 w_774_654# vdd 0.008451f
C712 p1 b1 0.022716f
C713 p3 w_726_513# 4.5e-19
C714 p2p1g0 vdd 0.439883f
C715 p1g0 w_440_301# 0.004305f
C716 p2g1 gnd 0.215208f
C717 p1g0 a_617_318# 4.37e-21
C718 a_453_311# p1p0c0 0.060798f
C719 w_329_n250# a2 0.007896f
C720 vdd w_620_464# 0.008451f
C721 a_302_n114# vdd 0.019283f
C722 b1 gnd 0.035378f
C723 w_879_518# vdd 0.013167f
C724 a_731_417# w_725_444# 0.008113f
C725 a_440_412# a_397_472# 0.41238f
C726 vdd w_505_625# 0.008451f
C727 a_771_282# cin 0.68509f
C728 w_238_456# a_218_418# 0.026794f
C729 b0 a_302_20# 0.685117f
C730 a_597_73# a_673_36# 0.060798f
C731 p0 a_445_147# 2.81e-20
C732 cin a_816_233# 0.002154f
C733 vdd w_347_461# 0.008451f
C734 p3p2p1g0 w_878_485# 0.011197f
C735 p2p1p0c0 a_693_378# 0.040556f
C736 w_581_n75# a_561_n113# 0.026794f
C737 w_657_n70# a_670_n102# 0.013216f
C738 w_584_63# p0 0.00465f
C739 a_445_140# w_439_167# 0.008113f
C740 w_611_272# a_617_278# 0.017071f
C741 w_676_271# a_600_239# 0.027289f
C742 w_758_272# a_771_282# 0.015055f
C743 a_600_239# gnd 0.829424f
C744 a_324_88# p0 0.0179f
C745 c1 a_597_73# 2.15e-19
C746 cin a_496_251# 0.014005f
C747 p0 a_304_190# 0.001371f
C748 g3 g1 0.023266f
C749 a_534_474# p2g1 9.1e-19
C750 w_548_n81# a1 0.02809f
C751 a_594_556# p2 0.023173f
C752 a_797_547# p3 0.013746f
C753 w_367_323# vdd 0.008493f
C754 a_381_614# w_472_604# 0.027163f
C755 g2 gnd 0.829522f
C756 p1 p0 0.070301f
C757 w_291_n117# vdd 0.008507f
C758 p3 a_688_664# 0.002444f
C759 w_611_305# p1g0 0.036784f
C760 p2 cin 0.005346f
C761 c4 gnd 0.20619f
C762 a_453_311# vdd 1.32165f
C763 b1 a_561_n113# 0.00343f
C764 a_269_20# gnd 0.248155f
C765 w_797_280# c2 0.003455f
C766 a_673_36# vdd 0.441416f
C767 a_534_474# w_521_464# 0.017642f
C768 gnd a_738_234# 0.206673f
C769 vdd a_380_153# 0.441416f
C770 a_302_20# w_367_22# 0.015055f
C771 g1 p2 0.146371f
C772 g2 b3 3.99e-19
C773 w_795_n349# p3 0.028034f
C774 a_518_635# vdd 1.76176f
C775 p0 gnd 0.67177f
C776 c1 vdd 0.439883f
C777 a_440_393# p1 0.013746f
C778 a_610_395# p0 0.019134f
C779 c1 c3 2.14e-19
C780 g3 p3p2g1 0.010274f
C781 a_594_556# a_594_575# 0.41238f
C782 a_884_498# p3g2 3.63e-19
C783 g2 a_206_556# 0.008991f
C784 a_594_n65# a1 0.001371f
C785 a_327_429# w_314_461# 0.013216f
C786 w_795_n349# a_808_n381# 0.013216f
C787 p3 a3 0.413834f
C788 c3 w_828_n343# 0.016729f
C789 w_834_277# vdd 0.008507f
C790 w_367_185# cin 0.00869f
C791 w_834_277# c3 3.18e-20
C792 a_440_393# gnd 0.41238f
C793 w_807_654# a_688_664# 0.027639f
C794 w_401_n240# p2 0.003504f
C795 w_400_n106# b1 0.015139f
C796 w_291_n117# a_302_n114# 0.027261f
C797 w_291_318# g0 0.008451f
C798 a_797_566# p3g2 0.004452f
C799 p1g0 g0 0.015977f
C800 p3g2 p1 0.057343f
C801 p3p2p1g0 p3 0.010267f
C802 p3p2g1 p2 0.017215f
C803 p2 a2 0.49284f
C804 vdd w_551_n357# 0.0086f
C805 a_564_n389# w_584_n351# 0.026794f
C806 a_673_n378# w_660_n346# 0.013216f
C807 a_325_n314# gnd 0.206673f
C808 a_564_n389# vdd 0.439891f
C809 w_258_17# vdd 0.008451f
C810 a_445_140# a_445_147# 0.453641f
C811 w_548_n81# p1 0.002922f
C812 p1 a_798_n113# 0.060798f
C813 p0 a_534_474# 0.005763f
C814 p2 p2g1 0.004909f
C815 b3 w_329_n384# 0.027716f
C816 b3 a_325_n314# 0.02927f
C817 p3p2p1p0c0 vdd 0.448649f
C818 p3g2 gnd 0.298314f
C819 a_518_635# w_505_625# 0.017642f
C820 a_883_429# a_883_389# 0.41238f
C821 p3p2p1g0 a_825_350# 0.040556f
C822 vdd a_325_n180# 0.439883f
C823 a_617_318# a_617_278# 0.41238f
C824 s2 a_873_n248# 0.20619f
C825 w_690_n70# vdd 0.008451f
C826 w_741_654# vdd 0.008451f
C827 p2 w_521_464# 0.026794f
C828 g1 a_670_n102# 0.060798f
C829 w_551_n219# a_564_n251# 0.013216f
C830 g1 a_397_472# 0.007928f
C831 p1 a1 0.008941f
C832 a_798_n113# gnd 0.206673f
C833 p1g0 w_400_323# 0.013216f
C834 a_218_418# gnd 0.20619f
C835 p2 w_401_604# 0.026996f
C836 p3p2g1 a_594_575# 7.98e-19
C837 a_731_417# a_693_378# 0.453641f
C838 p1g0 p1p0c0 0.011688f
C839 g1 w_417_462# 2.78e-19
C840 a_325_n180# a_329_n171# 0.14502f
C841 b2 a_564_n251# 0.002958f
C842 a_771_282# a_738_234# 0.286223f
C843 p1 a_594_n65# 0.004757f
C844 vdd w_587_464# 0.008451f
C845 a_738_234# a_816_233# 0.14502f
C846 a_269_n114# vdd 0.441416f
C847 a1 gnd 1.537765f
C848 w_726_513# vdd 0.013119f
C849 g3 g2 0.005441f
C850 a_440_412# g0 0.014522f
C851 p0 w_473_301# 0.026996f
C852 w_504_133# g0 0.011197f
C853 w_857_n67# s1 0.007992f
C854 vdd w_472_604# 0.008451f
C855 a_771_282# p0 0.413834f
C856 w_205_450# a_218_418# 0.013216f
C857 cin pocin 0.002387f
C858 a0 a_302_20# 0.413834f
C859 vdd w_314_461# 0.008507f
C860 a_594_n65# gnd 0.701773f
C861 p3p2p1p0c0 w_879_518# 0.015324f
C862 w_790_410# a_693_378# 0.027289f
C863 p3p2g1 w_878_485# 6.13e-19
C864 p2g1 a_693_378# 0.244568f
C865 p2p1p0c0 a_731_457# 4.37e-21
C866 g1 a_617_318# 0.010567f
C867 w_548_n81# a_561_n113# 0.013216f
C868 g2 p2 0.073455f
C869 w_551_57# p0 0.00465f
C870 w_611_272# a_600_239# 0.013329f
C871 w_611_305# a_617_278# 0.008113f
C872 a_847_245# gnd 0.248155f
C873 b0 p0 0.023585f
C874 p0 a_496_251# 0.013746f
C875 cin c2 0.003312f
C876 gnd a_445_147# 0.575941f
C877 a_251_466# g1 0.770057f
C878 a_397_472# p2g1 0.009943f
C879 a_797_566# p1 0.013746f
C880 a_594_556# p3 0.016756f
C881 a_424_554# p2 0.023081f
C882 w_291_318# vdd 6.13e-19
C883 a_381_614# w_434_604# 0.027639f
C884 p3g2 w_335_599# 0.013277f
C885 g1 c2 0.014621f
C886 w_258_n117# vdd 0.008451f
C887 p3 cin 0.00353f
C888 p2 p0 0.023721f
C889 a_380_291# gnd 0.248155f
C890 p1g0 vdd 0.451968f
C891 p2g1 w_417_462# 8.35e-22
C892 a_269_n114# a_302_n114# 0.060798f
C893 a_324_88# gnd 0.206673f
C894 a_324_n46# a_328_n37# 0.14502f
C895 a1 a_561_n113# 0.060856f
C896 w_758_272# c2 0.003448f
C897 gnd a_304_190# 0.701773f
C898 a_302_20# w_328_18# 0.007992f
C899 w_439_134# pocin 1.21e-19
C900 g1 p3 0.65866f
C901 p1 gnd 0.329008f
C902 a_688_664# vdd 2.20188f
C903 a_594_n65# a_561_n113# 0.003752f
C904 a_440_393# p2 0.013746f
C905 a_610_395# p1 0.013746f
C906 w_611_305# g1 0.002086f
C907 a_731_492# a_731_457# 0.41238f
C908 g2 a_693_378# 1.39e-20
C909 a_239_604# w_226_594# 0.019526f
C910 g3 p3g2 0.013858f
C911 p3 w_368_n380# 0.015055f
C912 w_795_n349# vdd 0.008518f
C913 p3 a_329_n305# 0.20619f
C914 w_797_280# vdd 0.001288f
C915 a_797_585# cin 2.05e-21
C916 a_797_604# a_688_664# 0.41238f
C917 w_797_280# c3 0.012687f
C918 s3 a_886_n382# 0.20619f
C919 w_291_180# cin 0.008451f
C920 w_368_n246# p2 0.018553f
C921 w_774_654# a_688_664# 0.027639f
C922 w_807_654# cin 0.026794f
C923 w_367_n112# b1 0.01395f
C924 a_731_492# w_725_479# 0.01128f
C925 w_291_n117# a_269_n114# 0.013216f
C926 w_400_n106# a1 0.028034f
C927 w_693_68# g0 0.01325f
C928 a_271_280# g0 0.001372f
C929 s1 c2 0.002762f
C930 p0 a_693_378# 6.43e-21
C931 a_564_n389# w_551_n357# 0.013216f
C932 p3p2g1 p3 0.017448f
C933 p3g2 p2 0.026294f
C934 vdd w_401_n374# 0.008451f
C935 w_660_n346# a_597_n341# 0.026907f
C936 a_673_n378# vdd 0.441416f
C937 b3 gnd 0.034146f
C938 vdd a3 0.20154f
C939 w_504_133# vdd 0.008451f
C940 w_675_654# p3 0.026794f
C941 w_551_n219# vdd 0.008518f
C942 p1 a_561_n113# 0.002494f
C943 g1 a_381_614# 0.059029f
C944 p2 a_218_418# 0.061185f
C945 p1 a_534_474# 0.015195f
C946 cin g0 0.016039f
C947 vdd w_226_594# 6.13e-19
C948 p3p2p1g0 vdd 0.447889f
C949 a_206_556# gnd 0.20619f
C950 w_854_n201# s2 0.007992f
C951 vdd b2 2.33e-19
C952 p1p0c0 a_617_278# 0.019123f
C953 a_771_282# a_847_245# 0.060798f
C954 p3p2g1 a_825_350# 0.001345f
C955 a_795_n247# a_873_n248# 0.14502f
C956 w_708_654# vdd 0.008451f
C957 w_657_n70# vdd 0.008507f
C958 g1 g0 6.14e-19
C959 a_561_n113# gnd 0.20619f
C960 p3p2p1g0 a_797_604# 0.043431f
C961 p3p2g1 a_797_585# 0.049949f
C962 w_584_n213# b2 0.008451f
C963 p2p1p0c0 vdd 0.439883f
C964 a_534_474# gnd 0.042086f
C965 p3g2 a_594_575# 0.042464f
C966 g3 a_847_245# 0.015251f
C967 a_304_328# g0 0.753587f
C968 a_731_417# a_731_457# 0.41238f
C969 p1g0 a_453_311# 0.010005f
C970 g1 w_384_462# 0.011399f
C971 a2 a_564_n251# 0.060856f
C972 b2 a_329_n171# 0.001802f
C973 a_600_239# c2 0.060798f
C974 vdd w_554_464# 0.008451f
C975 g1 a_327_429# 0.009049f
C976 a_324_n46# vdd 0.439891f
C977 p3p2p1p0c0 w_877_416# 0.018361f
C978 w_658_464# vdd 0.008451f
C979 a_381_614# p3p2g1 0.060798f
C980 a_315_567# p3g2 0.060798f
C981 p3p2p1p0c0 a_883_464# 0.005542f
C982 w_818_n75# s1 0.015055f
C983 w_439_134# g0 0.051057f
C984 w_400_n106# p1 3.76e-36
C985 vdd w_434_604# 0.008451f
C986 p1p0c0 cin 0.013387f
C987 b0 w_584_63# 0.008938f
C988 cin a_271_142# 0.001372f
C989 p0 pocin 5.46e-21
C990 b0 a_324_88# 0.02927f
C991 c2 a_738_234# 0.003282f
C992 a_886_n382# 0 0.016528f **FLOATING
C993 gnd 0 15.648485f **FLOATING
C994 s3 0 0.473154f **FLOATING
C995 a_808_n381# 0 0.526842f **FLOATING
C996 vdd 0 26.089828f **FLOATING
C997 a_564_n389# 0 0.477455f **FLOATING
C998 a_673_n378# 0 0.382299f **FLOATING
C999 a_329_n305# 0 0.016528f **FLOATING
C1000 a_325_n314# 0 0.526842f **FLOATING
C1001 b3 0 6.62907f **FLOATING
C1002 a3 0 2.45012f **FLOATING
C1003 a_597_n341# 0 0.771781f **FLOATING
C1004 a_873_n248# 0 0.016528f **FLOATING
C1005 s2 0 0.462937f **FLOATING
C1006 a_795_n247# 0 0.526842f **FLOATING
C1007 a_564_n251# 0 0.477455f **FLOATING
C1008 a_329_n171# 0 0.016528f **FLOATING
C1009 a_325_n180# 0 0.526842f **FLOATING
C1010 b2 0 6.55321f **FLOATING
C1011 a2 0 2.34823f **FLOATING
C1012 a_876_n114# 0 0.016528f **FLOATING
C1013 s1 0 0.462937f **FLOATING
C1014 a_798_n113# 0 0.526842f **FLOATING
C1015 a_561_n113# 0 0.477455f **FLOATING
C1016 a_670_n102# 0 0.382299f **FLOATING
C1017 a_328_n37# 0 0.016528f **FLOATING
C1018 a_302_n114# 0 0.662497f **FLOATING
C1019 a_269_n114# 0 0.382299f **FLOATING
C1020 a_324_n46# 0 0.526842f **FLOATING
C1021 b1 0 5.67427f **FLOATING
C1022 a1 0 2.37347f **FLOATING
C1023 a_594_n65# 0 0.771781f **FLOATING
C1024 a_564_25# 0 0.477455f **FLOATING
C1025 a_673_36# 0 0.382299f **FLOATING
C1026 a_328_97# 0 0.016528f **FLOATING
C1027 a_302_20# 0 0.662497f **FLOATING
C1028 a_269_20# 0 0.382299f **FLOATING
C1029 a_324_88# 0 0.526842f **FLOATING
C1030 b0 0 6.55446f **FLOATING
C1031 a0 0 2.49553f **FLOATING
C1032 a_597_73# 0 0.804448f **FLOATING
C1033 c1 0 2.24107f **FLOATING
C1034 a_445_140# 0 0.179875f **FLOATING
C1035 a_445_147# 0 1.02677f **FLOATING
C1036 a_816_233# 0 0.016528f **FLOATING
C1037 pocin 0 0.600283f **FLOATING
C1038 a_271_142# 0 0.477455f **FLOATING
C1039 a_380_153# 0 0.382299f **FLOATING
C1040 a_496_232# 0 0.040245f **FLOATING
C1041 s0 0 0.145867f **FLOATING
C1042 a_738_234# 0 0.526842f **FLOATING
C1043 a_304_190# 0 0.771781f **FLOATING
C1044 a_496_251# 0 0.040245f **FLOATING
C1045 c2 0 2.27948f **FLOATING
C1046 a_617_278# 0 0.206277f **FLOATING
C1047 a_600_239# 0 1.28245f **FLOATING
C1048 a_847_245# 0 0.382299f **FLOATING
C1049 a_771_282# 0 0.662497f **FLOATING
C1050 a_617_318# 0 0.150155f **FLOATING
C1051 p1p0c0 0 0.596493f **FLOATING
C1052 a_453_311# 0 1.70512f **FLOATING
C1053 p1g0 0 1.48359f **FLOATING
C1054 a_271_280# 0 0.477455f **FLOATING
C1055 c4 0 0.15567f **FLOATING
C1056 a_380_291# 0 0.382299f **FLOATING
C1057 a_610_377# 0 0.036687f **FLOATING
C1058 a_304_328# 0 0.771914f **FLOATING
C1059 a_440_393# 0 0.040245f **FLOATING
C1060 a_610_395# 0 0.040245f **FLOATING
C1061 a_883_389# 0 0.206277f **FLOATING
C1062 a_825_350# 0 1.81544f **FLOATING
C1063 c3 0 2.7802f **FLOATING
C1064 a_610_414# 0 0.040245f **FLOATING
C1065 a_440_412# 0 0.040245f **FLOATING
C1066 a_731_417# 0 0.206277f **FLOATING
C1067 a_883_429# 0 0.150155f **FLOATING
C1068 a_693_378# 0 1.54889f **FLOATING
C1069 a_731_457# 0 0.150155f **FLOATING
C1070 p2p1g0 0 0.681984f **FLOATING
C1071 a_883_464# 0 0.148414f **FLOATING
C1072 p2p1p0c0 0 1.73079f **FLOATING
C1073 p2g1 0 0.842448f **FLOATING
C1074 a_218_418# 0 0.477455f **FLOATING
C1075 a_534_474# 0 2.14225f **FLOATING
C1076 a_397_472# 0 1.70506f **FLOATING
C1077 g0 0 11.810905f **FLOATING
C1078 a_327_429# 0 0.382299f **FLOATING
C1079 a_731_492# 0 0.148414f **FLOATING
C1080 g2 0 17.347467f **FLOATING
C1081 a_884_498# 0 0.144831f **FLOATING
C1082 g3 0 6.01254f **FLOATING
C1083 a_251_466# 0 0.770807f **FLOATING
C1084 a_424_535# 0 0.040245f **FLOATING
C1085 a_594_537# 0 0.040245f **FLOATING
C1086 a_797_547# 0 0.040245f **FLOATING
C1087 a_594_556# 0 0.040245f **FLOATING
C1088 a_424_554# 0 0.040245f **FLOATING
C1089 a_797_566# 0 0.040245f **FLOATING
C1090 a_594_575# 0 0.040245f **FLOATING
C1091 a_797_585# 0 0.040245f **FLOATING
C1092 a_797_604# 0 0.040245f **FLOATING
C1093 p3p2p1p0c0 0 4.14703f **FLOATING
C1094 p3p2p1g0 0 6.28184f **FLOATING
C1095 p3p2g1 0 4.7141f **FLOATING
C1096 p3g2 0 5.75063f **FLOATING
C1097 a_206_556# 0 0.477455f **FLOATING
C1098 a_315_567# 0 0.382299f **FLOATING
C1099 a_381_614# 0 1.70511f **FLOATING
C1100 g1 0 21.5435f **FLOATING
C1101 a_239_604# 0 0.804448f **FLOATING
C1102 a_518_635# 0 2.1423f **FLOATING
C1103 a_688_664# 0 2.57948f **FLOATING
C1104 cin 0 4.56014f **FLOATING
C1105 p0 0 7.29675f **FLOATING
C1106 p1 0 13.9001f **FLOATING
C1107 p2 0 13.4629f **FLOATING
C1108 p3 0 14.903701f **FLOATING
C1109 w_867_n335# 0 1.25349f **FLOATING
C1110 w_828_n343# 0 1.34991f **FLOATING
C1111 w_795_n349# 0 1.34991f **FLOATING
C1112 w_693_n346# 0 1.34991f **FLOATING
C1113 w_660_n346# 0 1.34991f **FLOATING
C1114 w_584_n351# 0 1.34991f **FLOATING
C1115 w_551_n357# 0 1.34991f **FLOATING
C1116 w_401_n374# 0 1.34991f **FLOATING
C1117 w_368_n380# 0 1.34991f **FLOATING
C1118 w_329_n384# 0 1.25349f **FLOATING
C1119 w_854_n201# 0 1.25349f **FLOATING
C1120 w_815_n209# 0 1.34991f **FLOATING
C1121 w_782_n215# 0 1.34991f **FLOATING
C1122 w_584_n213# 0 1.34991f **FLOATING
C1123 w_551_n219# 0 1.34991f **FLOATING
C1124 w_401_n240# 0 1.34991f **FLOATING
C1125 w_368_n246# 0 1.34991f **FLOATING
C1126 w_329_n250# 0 1.25349f **FLOATING
C1127 w_857_n67# 0 1.25349f **FLOATING
C1128 w_818_n75# 0 1.34991f **FLOATING
C1129 w_785_n81# 0 1.34991f **FLOATING
C1130 w_690_n70# 0 1.34991f **FLOATING
C1131 w_657_n70# 0 1.34991f **FLOATING
C1132 w_581_n75# 0 1.34991f **FLOATING
C1133 w_548_n81# 0 1.34991f **FLOATING
C1134 w_400_n106# 0 1.34991f **FLOATING
C1135 w_367_n112# 0 1.34991f **FLOATING
C1136 w_328_n116# 0 1.25349f **FLOATING
C1137 w_291_n117# 0 1.34991f **FLOATING
C1138 w_258_n117# 0 1.34991f **FLOATING
C1139 w_693_68# 0 1.34991f **FLOATING
C1140 w_660_68# 0 1.34991f **FLOATING
C1141 w_584_63# 0 1.34991f **FLOATING
C1142 w_551_57# 0 1.34991f **FLOATING
C1143 w_400_28# 0 1.34991f **FLOATING
C1144 w_367_22# 0 1.34991f **FLOATING
C1145 w_328_18# 0 1.25349f **FLOATING
C1146 w_291_17# 0 1.34991f **FLOATING
C1147 w_258_17# 0 1.34991f **FLOATING
C1148 w_504_133# 0 1.34991f **FLOATING
C1149 w_439_134# 0 1.34991f **FLOATING
C1150 w_439_167# 0 1.34991f **FLOATING
C1151 w_400_185# 0 1.34991f **FLOATING
C1152 w_367_185# 0 1.34991f **FLOATING
C1153 w_291_180# 0 1.34991f **FLOATING
C1154 w_258_174# 0 1.34991f **FLOATING
C1155 w_867_277# 0 1.34991f **FLOATING
C1156 w_834_277# 0 1.34991f **FLOATING
C1157 w_797_280# 0 1.25349f **FLOATING
C1158 w_758_272# 0 1.34991f **FLOATING
C1159 w_725_266# 0 1.34991f **FLOATING
C1160 w_676_271# 0 1.34991f **FLOATING
C1161 w_611_272# 0 1.34991f **FLOATING
C1162 w_611_305# 0 1.34991f **FLOATING
C1163 w_611_340# 0 1.34991f **FLOATING
C1164 w_544_301# 0 1.34991f **FLOATING
C1165 w_506_301# 0 1.34991f **FLOATING
C1166 w_473_301# 0 1.34991f **FLOATING
C1167 w_440_301# 0 1.34991f **FLOATING
C1168 w_400_323# 0 1.34991f **FLOATING
C1169 w_367_323# 0 1.34991f **FLOATING
C1170 w_291_318# 0 1.34991f **FLOATING
C1171 w_258_312# 0 1.34991f **FLOATING
C1172 w_942_382# 0 1.34991f **FLOATING
C1173 w_877_383# 0 1.34991f **FLOATING
C1174 w_877_416# 0 1.34991f **FLOATING
C1175 w_877_451# 0 1.34991f **FLOATING
C1176 w_790_410# 0 1.34991f **FLOATING
C1177 w_725_411# 0 1.34991f **FLOATING
C1178 w_725_444# 0 1.34991f **FLOATING
C1179 w_878_485# 0 1.34991f **FLOATING
C1180 w_725_479# 0 1.34991f **FLOATING
C1181 w_879_518# 0 1.34991f **FLOATING
C1182 w_726_513# 0 1.34991f **FLOATING
C1183 w_658_464# 0 1.34991f **FLOATING
C1184 w_620_464# 0 1.34991f **FLOATING
C1185 w_587_464# 0 1.34991f **FLOATING
C1186 w_554_464# 0 1.34991f **FLOATING
C1187 w_521_464# 0 1.34991f **FLOATING
C1188 w_488_462# 0 1.34991f **FLOATING
C1189 w_450_462# 0 1.34991f **FLOATING
C1190 w_417_462# 0 1.34991f **FLOATING
C1191 w_384_462# 0 1.34991f **FLOATING
C1192 w_347_461# 0 1.34991f **FLOATING
C1193 w_314_461# 0 1.34991f **FLOATING
C1194 w_238_456# 0 1.34991f **FLOATING
C1195 w_205_450# 0 1.34991f **FLOATING
C1196 w_845_654# 0 1.34991f **FLOATING
C1197 w_807_654# 0 1.34991f **FLOATING
C1198 w_774_654# 0 1.34991f **FLOATING
C1199 w_741_654# 0 1.34991f **FLOATING
C1200 w_708_654# 0 1.34991f **FLOATING
C1201 w_675_654# 0 1.34991f **FLOATING
C1202 w_642_625# 0 1.34991f **FLOATING
C1203 w_604_625# 0 1.34991f **FLOATING
C1204 w_571_625# 0 1.34991f **FLOATING
C1205 w_538_625# 0 1.34991f **FLOATING
C1206 w_505_625# 0 1.34991f **FLOATING
C1207 w_472_604# 0 1.34991f **FLOATING
C1208 w_434_604# 0 1.34991f **FLOATING
C1209 w_401_604# 0 1.34991f **FLOATING
C1210 w_368_604# 0 1.34991f **FLOATING
C1211 w_335_599# 0 1.34991f **FLOATING
C1212 w_302_599# 0 1.34991f **FLOATING
C1213 w_226_594# 0 1.34991f **FLOATING
C1214 w_193_588# 0 1.34991f **FLOATING
