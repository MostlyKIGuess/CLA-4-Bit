magic
tech scmos
timestamp 1731076245
<< nwell >>
rect 569 57 593 113
rect 602 63 626 119
rect 678 68 702 124
rect 711 68 735 124
rect 566 -81 590 -25
rect 599 -75 623 -19
rect 675 -70 699 -14
rect 708 -70 732 -14
rect 569 -219 593 -163
rect 602 -213 626 -157
rect 678 -208 702 -152
rect 711 -208 735 -152
rect 569 -357 593 -301
rect 602 -351 626 -295
rect 678 -346 702 -290
rect 711 -346 735 -290
<< ntransistor >>
rect 628 136 648 138
rect 628 50 648 52
rect 580 25 582 45
rect 689 36 691 56
rect 722 36 724 56
rect 625 -2 645 0
rect 625 -88 645 -86
rect 577 -113 579 -93
rect 686 -102 688 -82
rect 719 -102 721 -82
rect 628 -140 648 -138
rect 628 -226 648 -224
rect 580 -251 582 -231
rect 689 -240 691 -220
rect 722 -240 724 -220
rect 628 -278 648 -276
rect 628 -364 648 -362
rect 580 -389 582 -369
rect 689 -378 691 -358
rect 722 -378 724 -358
<< ptransistor >>
rect 580 67 582 107
rect 613 73 615 113
rect 689 78 691 118
rect 722 78 724 118
rect 577 -71 579 -31
rect 610 -65 612 -25
rect 686 -60 688 -20
rect 719 -60 721 -20
rect 580 -209 582 -169
rect 613 -203 615 -163
rect 689 -198 691 -158
rect 722 -198 724 -158
rect 580 -347 582 -307
rect 613 -341 615 -301
rect 689 -336 691 -296
rect 722 -336 724 -296
<< ndiffusion >>
rect 628 138 648 139
rect 628 135 648 136
rect 628 52 648 53
rect 628 49 648 50
rect 579 25 580 45
rect 582 25 583 45
rect 688 36 689 56
rect 691 36 692 56
rect 721 36 722 56
rect 724 36 725 56
rect 625 0 645 1
rect 625 -3 645 -2
rect 625 -86 645 -85
rect 625 -89 645 -88
rect 576 -113 577 -93
rect 579 -113 580 -93
rect 685 -102 686 -82
rect 688 -102 689 -82
rect 718 -102 719 -82
rect 721 -102 722 -82
rect 628 -138 648 -137
rect 628 -141 648 -140
rect 628 -224 648 -223
rect 628 -227 648 -226
rect 579 -251 580 -231
rect 582 -251 583 -231
rect 688 -240 689 -220
rect 691 -240 692 -220
rect 721 -240 722 -220
rect 724 -240 725 -220
rect 628 -276 648 -275
rect 628 -279 648 -278
rect 628 -362 648 -361
rect 628 -365 648 -364
rect 579 -389 580 -369
rect 582 -389 583 -369
rect 688 -378 689 -358
rect 691 -378 692 -358
rect 721 -378 722 -358
rect 724 -378 725 -358
<< pdiffusion >>
rect 579 67 580 107
rect 582 67 583 107
rect 612 73 613 113
rect 615 73 616 113
rect 688 78 689 118
rect 691 78 692 118
rect 721 78 722 118
rect 724 78 725 118
rect 576 -71 577 -31
rect 579 -71 580 -31
rect 609 -65 610 -25
rect 612 -65 613 -25
rect 685 -60 686 -20
rect 688 -60 689 -20
rect 718 -60 719 -20
rect 721 -60 722 -20
rect 579 -209 580 -169
rect 582 -209 583 -169
rect 612 -203 613 -163
rect 615 -203 616 -163
rect 688 -198 689 -158
rect 691 -198 692 -158
rect 721 -198 722 -158
rect 724 -198 725 -158
rect 579 -347 580 -307
rect 582 -347 583 -307
rect 612 -341 613 -301
rect 615 -341 616 -301
rect 688 -336 689 -296
rect 691 -336 692 -296
rect 721 -336 722 -296
rect 724 -336 725 -296
<< ndcontact >>
rect 628 139 648 143
rect 628 131 648 135
rect 628 53 648 57
rect 628 45 648 49
rect 575 25 579 45
rect 583 25 587 45
rect 684 36 688 56
rect 692 36 696 56
rect 717 36 721 56
rect 725 36 729 56
rect 625 1 645 5
rect 625 -7 645 -3
rect 625 -85 645 -81
rect 625 -93 645 -89
rect 572 -113 576 -93
rect 580 -113 584 -93
rect 681 -102 685 -82
rect 689 -102 693 -82
rect 714 -102 718 -82
rect 722 -102 726 -82
rect 628 -137 648 -133
rect 628 -145 648 -141
rect 628 -223 648 -219
rect 628 -231 648 -227
rect 575 -251 579 -231
rect 583 -251 587 -231
rect 684 -240 688 -220
rect 692 -240 696 -220
rect 717 -240 721 -220
rect 725 -240 729 -220
rect 628 -275 648 -271
rect 628 -283 648 -279
rect 628 -361 648 -357
rect 628 -369 648 -365
rect 575 -389 579 -369
rect 583 -389 587 -369
rect 684 -378 688 -358
rect 692 -378 696 -358
rect 717 -378 721 -358
rect 725 -378 729 -358
<< pdcontact >>
rect 575 67 579 107
rect 583 67 587 107
rect 608 73 612 113
rect 616 73 620 113
rect 684 78 688 118
rect 692 78 696 118
rect 717 78 721 118
rect 725 78 729 118
rect 572 -71 576 -31
rect 580 -71 584 -31
rect 605 -65 609 -25
rect 613 -65 617 -25
rect 681 -60 685 -20
rect 689 -60 693 -20
rect 714 -60 718 -20
rect 722 -60 726 -20
rect 575 -209 579 -169
rect 583 -209 587 -169
rect 608 -203 612 -163
rect 616 -203 620 -163
rect 684 -198 688 -158
rect 692 -198 696 -158
rect 717 -198 721 -158
rect 725 -198 729 -158
rect 575 -347 579 -307
rect 583 -347 587 -307
rect 608 -341 612 -301
rect 616 -341 620 -301
rect 684 -336 688 -296
rect 692 -336 696 -296
rect 717 -336 721 -296
rect 725 -336 729 -296
<< polysilicon >>
rect 625 136 628 138
rect 648 136 651 138
rect 689 118 691 121
rect 722 118 724 121
rect 613 113 615 116
rect 580 107 582 110
rect 580 45 582 67
rect 613 61 615 73
rect 689 56 691 78
rect 722 56 724 78
rect 620 50 628 52
rect 648 50 651 52
rect 689 33 691 36
rect 722 33 724 36
rect 580 22 582 25
rect 622 -2 625 0
rect 645 -2 648 0
rect 686 -20 688 -17
rect 719 -20 721 -17
rect 610 -25 612 -22
rect 577 -31 579 -28
rect 577 -93 579 -71
rect 610 -77 612 -65
rect 686 -82 688 -60
rect 719 -82 721 -60
rect 617 -88 625 -86
rect 645 -88 648 -86
rect 686 -105 688 -102
rect 719 -105 721 -102
rect 577 -116 579 -113
rect 625 -140 628 -138
rect 648 -140 651 -138
rect 689 -158 691 -155
rect 722 -158 724 -155
rect 613 -163 615 -160
rect 580 -169 582 -166
rect 580 -231 582 -209
rect 613 -215 615 -203
rect 689 -220 691 -198
rect 722 -220 724 -198
rect 620 -226 628 -224
rect 648 -226 651 -224
rect 689 -243 691 -240
rect 722 -243 724 -240
rect 580 -254 582 -251
rect 625 -278 628 -276
rect 648 -278 651 -276
rect 689 -296 691 -293
rect 722 -296 724 -293
rect 613 -301 615 -298
rect 580 -307 582 -304
rect 580 -369 582 -347
rect 613 -353 615 -341
rect 689 -358 691 -336
rect 722 -358 724 -336
rect 620 -364 628 -362
rect 648 -364 651 -362
rect 689 -381 691 -378
rect 722 -381 724 -378
rect 580 -392 582 -389
<< polycontact >>
rect 621 135 625 139
rect 576 49 580 53
rect 612 57 616 61
rect 685 60 689 64
rect 718 60 722 64
rect 616 49 620 53
rect 618 -3 622 1
rect 573 -89 577 -85
rect 609 -81 613 -77
rect 682 -78 686 -74
rect 715 -78 719 -74
rect 613 -89 617 -85
rect 621 -141 625 -137
rect 576 -227 580 -223
rect 612 -219 616 -215
rect 685 -216 689 -212
rect 718 -216 722 -212
rect 616 -227 620 -223
rect 621 -279 625 -275
rect 576 -365 580 -361
rect 612 -357 616 -353
rect 685 -354 689 -350
rect 718 -354 722 -350
rect 616 -365 620 -361
<< metal1 >>
rect 648 139 661 143
rect 561 135 621 139
rect 561 53 566 135
rect 644 122 648 131
rect 569 113 593 120
rect 602 119 648 122
rect 608 113 612 119
rect 575 107 579 113
rect 583 53 587 67
rect 616 68 620 73
rect 655 68 661 139
rect 678 124 735 131
rect 684 118 688 124
rect 717 118 721 124
rect 616 65 661 68
rect 616 64 678 65
rect 692 64 696 78
rect 725 64 729 78
rect 612 53 616 57
rect 648 53 652 64
rect 658 60 685 64
rect 692 60 718 64
rect 725 60 737 64
rect 692 56 696 60
rect 725 56 729 60
rect 561 49 576 53
rect 583 49 616 53
rect 583 45 587 49
rect -90 20 -42 33
rect 470 25 518 38
rect -90 4 -42 17
rect 470 9 518 22
rect 575 16 579 25
rect 644 16 648 45
rect 684 16 688 36
rect 717 16 721 36
rect 569 8 736 16
rect 645 1 658 5
rect 558 -3 618 1
rect 558 -85 563 -3
rect 641 -16 645 -7
rect 566 -25 590 -18
rect 599 -19 645 -16
rect 605 -25 609 -19
rect 572 -31 576 -25
rect 580 -85 584 -71
rect 613 -70 617 -65
rect 652 -70 658 1
rect 675 -14 732 -7
rect 681 -20 685 -14
rect 714 -20 718 -14
rect 613 -73 658 -70
rect 613 -74 675 -73
rect 689 -74 693 -60
rect 722 -74 726 -60
rect 609 -85 613 -81
rect 645 -85 649 -74
rect 655 -78 682 -74
rect 689 -78 715 -74
rect 722 -78 734 -74
rect 689 -82 693 -78
rect 722 -82 726 -78
rect 558 -89 573 -85
rect 580 -89 613 -85
rect 580 -93 584 -89
rect -90 -117 -42 -104
rect 470 -112 518 -99
rect -90 -132 -42 -120
rect 470 -127 518 -115
rect 572 -122 576 -113
rect 641 -122 645 -93
rect 681 -122 685 -102
rect 714 -122 718 -102
rect 566 -130 733 -122
rect 648 -137 661 -133
rect 561 -141 621 -137
rect 561 -223 566 -141
rect 644 -154 648 -145
rect 569 -163 593 -156
rect 602 -157 648 -154
rect 608 -163 612 -157
rect 575 -169 579 -163
rect 583 -223 587 -209
rect 616 -208 620 -203
rect 655 -208 661 -137
rect 678 -152 735 -145
rect 684 -158 688 -152
rect 717 -158 721 -152
rect 616 -211 661 -208
rect 616 -212 678 -211
rect 692 -212 696 -198
rect 725 -212 729 -198
rect 612 -223 616 -219
rect 648 -223 652 -212
rect 658 -216 685 -212
rect 692 -216 718 -212
rect 725 -216 737 -212
rect 692 -220 696 -216
rect 725 -220 729 -216
rect 561 -227 576 -223
rect 583 -227 616 -223
rect 583 -231 587 -227
rect -90 -254 -42 -242
rect 470 -249 518 -237
rect -90 -270 -42 -257
rect 470 -265 518 -252
rect 575 -260 579 -251
rect 644 -260 648 -231
rect 684 -260 688 -240
rect 717 -260 721 -240
rect 569 -268 736 -260
rect 648 -275 661 -271
rect 561 -279 621 -275
rect 561 -361 566 -279
rect 644 -292 648 -283
rect 569 -301 593 -294
rect 602 -295 648 -292
rect 608 -301 612 -295
rect 575 -307 579 -301
rect 583 -361 587 -347
rect 616 -346 620 -341
rect 655 -346 661 -275
rect 678 -290 735 -283
rect 684 -296 688 -290
rect 717 -296 721 -290
rect 616 -349 661 -346
rect 616 -350 678 -349
rect 692 -350 696 -336
rect 725 -350 729 -336
rect 612 -361 616 -357
rect 648 -361 652 -350
rect 658 -354 685 -350
rect 692 -354 718 -350
rect 725 -354 737 -350
rect 692 -358 696 -354
rect 725 -358 729 -354
rect 561 -365 576 -361
rect 583 -365 616 -361
rect 583 -369 587 -365
rect -90 -395 -42 -382
rect 470 -390 518 -377
rect -90 -411 -42 -398
rect 470 -406 518 -393
rect 575 -398 579 -389
rect 644 -398 648 -369
rect 684 -398 688 -378
rect 717 -398 721 -378
rect 569 -406 736 -398
rect -90 -452 -42 -439
rect 470 -447 518 -434
<< metal2 >>
rect 584 124 678 131
rect 584 120 592 124
rect 73 16 78 115
rect 170 53 204 61
rect 633 21 638 120
rect 730 58 764 66
rect 507 16 638 21
rect -53 11 78 16
rect 581 -14 675 -7
rect 581 -18 589 -14
rect 68 -121 75 -24
rect 173 -85 204 -77
rect 628 -116 635 -19
rect 733 -80 764 -72
rect 504 -121 635 -116
rect -56 -126 75 -121
rect 584 -152 678 -145
rect 584 -156 592 -152
rect 77 -259 82 -161
rect 174 -223 208 -216
rect 637 -254 642 -156
rect 734 -218 768 -211
rect 512 -259 642 -254
rect -48 -264 82 -259
rect 584 -290 678 -283
rect 584 -294 592 -290
rect 75 -398 80 -300
rect 174 -361 209 -354
rect 635 -393 640 -295
rect 734 -356 769 -349
rect 511 -397 640 -393
rect -49 -402 80 -398
<< metal3 >>
rect -57 42 12 50
rect 503 47 572 55
rect -57 27 -52 42
rect 503 32 508 47
rect 506 -88 571 -83
rect -54 -93 11 -88
rect -54 -107 -47 -93
rect 506 -102 513 -88
rect -50 -234 14 -228
rect 510 -229 574 -223
rect -50 -245 -45 -234
rect 510 -240 515 -229
rect -53 -372 15 -366
rect 507 -367 575 -361
rect -53 -384 -46 -372
rect 507 -379 514 -367
<< pad >>
rect 678 124 686 131
rect 73 109 81 117
rect 584 113 592 120
rect 633 114 641 122
rect 170 53 178 61
rect 730 58 738 66
rect 12 42 20 50
rect 572 47 580 55
rect -58 25 -50 33
rect 502 30 510 38
rect -53 9 -45 17
rect 507 14 515 22
rect 675 -14 683 -7
rect 68 -28 75 -21
rect 581 -25 589 -18
rect 628 -23 635 -16
rect 170 -85 178 -77
rect 730 -80 738 -72
rect 10 -95 17 -88
rect 570 -90 577 -83
rect -56 -113 -46 -104
rect 504 -108 514 -99
rect -56 -129 -46 -120
rect 504 -124 514 -115
rect 678 -152 686 -145
rect 77 -166 84 -159
rect 584 -163 592 -156
rect 637 -161 644 -154
rect 174 -223 181 -216
rect 734 -218 741 -211
rect 13 -234 20 -227
rect 573 -229 580 -222
rect -52 -249 -45 -242
rect 508 -244 515 -237
rect -51 -264 -44 -257
rect 509 -259 516 -252
rect 678 -290 686 -283
rect 75 -304 82 -297
rect 584 -301 592 -294
rect 635 -299 642 -292
rect 174 -361 181 -354
rect 734 -356 741 -349
rect 13 -372 20 -365
rect 573 -367 580 -360
rect -53 -389 -46 -382
rect 507 -384 514 -377
rect -51 -405 -44 -398
rect 509 -400 516 -393
use and  and_0
timestamp 1731006496
transform 1 0 25 0 1 54
box -24 -51 152 84
use and  and_1
timestamp 1731006496
transform 1 0 22 0 1 -84
box -24 -51 152 84
use and  and_2
timestamp 1731006496
transform 1 0 25 0 1 -222
box -24 -51 152 84
use and  and_3
timestamp 1731006496
transform 1 0 25 0 1 -360
box -24 -51 152 84
<< labels >>
rlabel metal1 -71 27 -71 27 1 a0
rlabel metal1 -72 10 -72 10 1 a1
rlabel metal2 194 58 194 58 1 g0
rlabel metal1 -72 -110 -72 -110 1 a2
rlabel metal1 -72 -125 -72 -125 1 a3
rlabel metal2 193 -81 193 -81 1 g1
rlabel metal1 -71 -248 -71 -248 1 b0
rlabel metal1 -72 -263 -72 -263 1 b1
rlabel metal2 192 -220 192 -220 1 g2
rlabel metal1 -72 -448 -72 -448 1 c0
rlabel metal1 -67 -390 -67 -390 1 b2
rlabel metal1 -71 -402 -71 -402 1 b3
rlabel metal2 196 -357 196 -357 1 g3
rlabel metal1 489 32 489 32 1 a0
rlabel metal1 488 15 488 15 1 a1
rlabel metal2 754 63 754 63 1 g0
rlabel metal1 488 -105 488 -105 1 a2
rlabel metal1 488 -120 488 -120 1 a3
rlabel metal2 753 -76 753 -76 1 g1
rlabel metal1 489 -243 489 -243 1 b0
rlabel metal1 488 -258 488 -258 1 b1
rlabel metal2 752 -215 752 -215 1 g2
rlabel metal1 488 -443 488 -443 1 c0
rlabel metal1 493 -385 493 -385 1 b2
rlabel metal1 489 -397 489 -397 1 b3
rlabel metal2 756 -352 756 -352 1 g3
rlabel metal1 568 -365 574 -362 3 a
rlabel metal1 592 -365 597 -363 7 abar
rlabel metal1 580 -299 580 -299 5 vdd
rlabel metal1 609 -293 609 -293 1 b
rlabel metal1 705 -352 705 -352 1 ybar
rlabel metal1 732 -352 732 -352 7 y
rlabel metal1 689 -288 689 -288 5 vdd
rlabel metal1 722 -288 722 -288 5 vdd
rlabel metal1 657 -312 657 -312 1 y-d
rlabel metal1 575 -402 575 -402 1 gnd
rlabel metal1 568 -227 574 -224 3 a
rlabel metal1 592 -227 597 -225 7 abar
rlabel metal1 580 -161 580 -161 5 vdd
rlabel metal1 609 -155 609 -155 1 b
rlabel metal1 705 -214 705 -214 1 ybar
rlabel metal1 732 -214 732 -214 7 y
rlabel metal1 689 -150 689 -150 5 vdd
rlabel metal1 722 -150 722 -150 5 vdd
rlabel metal1 657 -174 657 -174 1 y-d
rlabel metal1 575 -264 575 -264 1 gnd
rlabel metal1 565 -89 571 -86 3 a
rlabel metal1 589 -89 594 -87 7 abar
rlabel metal1 577 -23 577 -23 5 vdd
rlabel metal1 606 -17 606 -17 1 b
rlabel metal1 702 -76 702 -76 1 ybar
rlabel metal1 729 -76 729 -76 7 y
rlabel metal1 686 -12 686 -12 5 vdd
rlabel metal1 719 -12 719 -12 5 vdd
rlabel metal1 654 -36 654 -36 1 y-d
rlabel metal1 572 -126 572 -126 1 gnd
rlabel metal1 568 49 574 52 3 a
rlabel metal1 592 49 597 51 7 abar
rlabel metal1 580 115 580 115 5 vdd
rlabel metal1 609 121 609 121 1 b
rlabel metal1 705 62 705 62 1 ybar
rlabel metal1 732 62 732 62 7 y
rlabel metal1 689 126 689 126 5 vdd
rlabel metal1 722 126 722 126 5 vdd
rlabel metal1 657 102 657 102 1 y-d
rlabel metal1 575 12 575 12 1 gnd
<< end >>
