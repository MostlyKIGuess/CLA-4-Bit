* SPICE3 file created from testing.ext - technology: scmos

.option scale=90n

M1000 a_594_537# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1001 a_239_604# p3 g2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_329_n305# a_325_n314# p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 a_218_418# p2 vdd w_205_450# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_825_350# g3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1005 a_600_239# p1p0c0 a_617_278# w_611_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 s1 p1 c1 w_818_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 c1 a_445_147# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1008 p3p2p1g0 a_518_635# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1009 a_693_378# p2g1 a_731_417# w_725_411# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_564_n251# a2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1011 a_600_239# p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 a_594_n65# a1 b1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 gnd a_269_20# p0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 a_594_556# p2 a_594_537# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 a_445_147# g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1016 a_594_575# p1 a_594_556# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1017 p2g1 a_327_429# vdd w_347_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1018 a_440_412# p1 a_440_393# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_564_n389# a3 vdd w_551_n357# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1020 p1p0c0 a_453_311# vdd w_544_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1021 a3 b3 p3 w_329_n384# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 a_518_635# p3 vdd w_505_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a_731_457# p2p1p0c0 a_731_417# w_725_444# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1024 a_808_n381# p3 vdd w_795_n349# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1025 b2 a2 p2 w_368_n246# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1026 p3p2g1 a_381_614# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 p2p1p0c0 a_534_474# vdd w_658_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1028 a_610_395# p1 a_610_377# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1029 a_329_n171# a_325_n180# p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 a_518_635# g0 a_594_575# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 s2 a_795_n247# a_873_n248# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 vdd a0 a_324_88# w_400_28# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1033 a_594_n65# a_561_n113# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1034 vdd a_302_20# a_269_20# w_291_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 a_325_n180# b2 p2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 a_825_350# p3p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1037 a_304_190# a_271_142# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1038 a_847_245# a_771_282# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1039 a_884_498# p3g2 a_883_464# w_878_485# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 a_731_492# p2p1g0 a_731_457# w_725_479# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1041 a_673_n378# a_597_n341# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 a_597_n341# a_564_n389# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1043 a_315_567# a_239_604# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 g0 a_673_36# vdd w_693_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 p3g2 a_315_567# vdd w_335_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 vdd g3 a_884_498# w_879_518# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1047 a_825_350# p3p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 pocin a_380_153# vdd w_400_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 vdd a_269_20# p0 w_258_17# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 a_218_418# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1051 a_380_153# a_304_190# vdd w_367_185# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 b1 a1 a_302_n114# w_367_n112# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_825_350# p3p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1054 a_271_280# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1055 p3p2p1g0 a_518_635# vdd w_642_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_239_604# a_206_556# g2 w_226_594# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 a_304_190# a_271_142# cin w_291_180# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 c3 a_693_378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 g3 a_673_n378# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 p2p1g0 a_397_472# vdd w_488_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_440_393# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_688_664# p0 vdd w_774_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 s2 p2 c2 w_815_n209# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1064 a_445_147# pocin gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 p2g1 a_327_429# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 a_600_239# p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1067 a_795_n247# p2 vdd w_782_n215# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_564_n251# a2 vdd w_551_n219# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_327_429# a_251_466# vdd w_314_461# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 a_688_664# cin vdd w_807_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1071 a_693_378# p2g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_251_466# p2 g1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 s1 c1 a_798_n113# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_798_n113# p1 vdd w_785_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_325_n314# b3 p3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 a_738_234# p0 vdd w_725_266# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1077 a_673_36# a_597_73# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1078 a_564_25# a0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1079 p3p2g1 a_381_614# vdd w_472_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1080 a_597_n341# a_564_n389# b3 w_584_n351# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1081 a_206_556# p3 vdd w_193_588# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_424_535# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1083 g2 a_564_n251# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1084 g1 a_670_n102# vdd w_690_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1085 s3 p3 c3 w_828_n343# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_610_377# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1087 s0 a_847_245# vdd w_867_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1088 vdd a2 a_325_n180# w_401_n240# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_670_n102# a_594_n65# vdd w_657_n70# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 c4 a_825_350# vdd w_942_382# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_670_n102# a_594_n65# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_424_554# p2 a_424_535# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 a_453_311# p0 vdd w_473_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1094 a_315_567# a_239_604# vdd w_302_599# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 p3p2p1p0c0 a_688_664# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_771_282# p0 cin w_758_272# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1097 s1 c1 p1 w_857_n67# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_271_142# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1099 a_534_474# cin vdd w_620_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_534_474# p0 vdd w_587_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_453_311# cin vdd w_506_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1102 a_271_280# p1 vdd w_258_312# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_561_n113# a1 vdd w_548_n81# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 a_381_614# g1 a_424_554# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_883_429# p3p2p1g0 a_883_389# w_877_416# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_693_378# p2p1g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 c1 a_445_147# vdd w_504_133# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_304_328# a_271_280# g0 w_291_318# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 a_825_350# p3g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1110 a_564_n389# a3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 s1 a_798_n113# a_876_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_688_664# p1 vdd w_741_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1113 a_797_604# p0 a_797_585# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 vdd a_269_n114# p1 w_258_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1115 p1g0 a_380_291# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_324_n46# b1 a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 a_327_429# a_251_466# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1118 a_693_378# p2p1p0c0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 a_380_291# a_304_328# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1120 c2 a_600_239# vdd w_676_271# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 b3 a3 p3 w_368_n380# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1122 a1 b1 a_302_n114# w_328_n116# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 a_328_n37# a_324_n46# a_302_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1124 a_328_97# a_324_88# a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 vdd a3 a_325_n314# w_401_n374# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1126 a_597_n341# a3 b3 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 p1p0c0 a_453_311# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1128 a_324_88# b0 a_302_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1129 a_688_664# cin a_797_604# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 vdd g2 a_731_492# w_726_513# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1131 a_883_464# p3p2g1 a_883_429# w_877_451# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_693_378# g2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_304_328# p1 g0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1134 g2 a_564_n251# b2 w_584_n213# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1135 a_597_73# a_564_25# b0 w_584_63# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1136 a_597_73# a0 b0 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1137 a_771_282# a_738_234# a_816_233# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1138 a_518_635# p1 vdd w_571_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_397_472# g0 vdd w_450_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_797_547# p3 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_496_251# p0 a_496_232# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 a_847_245# a_771_282# vdd w_834_277# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_597_73# a_564_25# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1147 a_239_604# a_206_556# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1148 a_797_566# p2 a_797_547# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1149 a_453_311# cin a_496_251# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1150 a_453_311# p1 vdd w_440_301# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 gnd a3 a_325_n314# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1152 a_534_474# p1 vdd w_554_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_304_328# a_271_280# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1154 a_445_147# g0 a_445_140# w_439_134# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 a_797_585# p1 a_797_566# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 gnd a_302_n114# a_269_n114# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_795_n247# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1158 gnd a_269_n114# p1 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1159 g0 a_673_36# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1160 a_381_614# g1 vdd w_434_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 s2 c2 a_795_n247# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_561_n113# a1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1163 pocin a_380_153# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_380_153# a_304_190# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1165 a_688_664# p3 vdd w_675_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1166 s3 a_808_n381# a_886_n382# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1167 a_673_n378# a_597_n341# vdd w_660_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 g2 a2 b2 Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 p1g0 a_380_291# vdd w_400_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1170 c2 a_600_239# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 g1 a_670_n102# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1172 a0 b0 a_302_20# w_328_18# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 a_380_291# a_304_328# vdd w_367_323# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_688_664# p2 vdd w_708_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1175 p2p1g0 a_397_472# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1176 gnd a2 a_325_n180# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 vdd pocin a_445_140# w_439_167# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1178 c3 a_693_378# vdd w_790_410# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_304_190# p0 cin Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1180 s3 c3 a_808_n381# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1181 a_251_466# a_218_418# g1 w_238_456# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1182 s3 c3 p3 w_867_n335# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 vdd a1 a_324_n46# w_400_n106# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1184 a_673_36# a_597_73# vdd w_660_68# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1185 a_397_472# g0 a_440_412# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 a_808_n381# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1187 a_798_n113# p1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_564_25# a0 vdd w_551_57# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 g3 a_673_n378# vdd w_693_n346# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# p2 vdd w_384_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 vdd a_302_n114# a_269_n114# w_291_n117# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1192 a_617_318# p1g0 a_617_278# w_611_305# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1193 a_771_282# cin p0 w_797_280# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 a_738_234# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1195 a_594_n65# a_561_n113# b1 w_581_n75# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_518_635# p2 vdd w_538_625# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 b0 a0 a_302_20# w_367_22# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_496_232# p1 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1199 a_397_472# p1 vdd w_417_462# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_206_556# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1201 p3p2p1p0c0 a_688_664# vdd w_845_654# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 a_610_414# p0 a_610_395# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_534_474# p2 vdd w_521_464# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_271_142# p0 vdd w_258_174# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1205 s0 a_847_245# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 vdd g1 a_617_318# w_611_340# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 c4 a_825_350# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1208 gnd a1 a_324_n46# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1209 gnd a0 a_324_88# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 gnd a_302_20# a_269_20# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1211 a_381_614# p2 vdd w_401_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1212 a2 b2 p2 w_329_n250# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 a_251_466# a_218_418# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 a_534_474# cin a_610_414# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1215 a_771_282# cin a_738_234# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 a_381_614# p3 vdd w_368_604# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1217 p3g2 a_315_567# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1218 a_600_239# g1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1219 s2 c2 p2 w_854_n201# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 a_304_328# a_271_280# 0.003752f
C1 w_834_277# a_847_245# 0.013216f
C2 w_725_266# c2 0.003448f
C3 p3 a_325_n314# 0.286223f
C4 gnd a_594_n65# 0.701773f
C5 p1 w_785_n81# 0.028309f
C6 p1 w_548_n81# 0.002922f
C7 gnd p3p2g1 0.234908f
C8 w_815_n209# c2 0.01623f
C9 p2 a_424_554# 0.023081f
C10 p1 a_797_566# 0.013746f
C11 cin a_600_239# 8.95e-19
C12 p1 c2 0.003604f
C13 a_440_412# gnd 1.91e-19
C14 gnd a_610_377# 0.41238f
C15 b2 w_329_n250# 0.027716f
C16 a2 w_368_n246# 0.028748f
C17 w_611_340# g1 0.039692f
C18 p1g0 a_453_311# 0.010005f
C19 p0 p2p1g0 0.009782f
C20 cin p2g1 0.013147f
C21 p0 w_660_68# 0.004686f
C22 vdd w_417_462# 0.008451f
C23 a_688_664# w_845_654# 0.027163f
C24 a_600_239# g1 1.39e-20
C25 w_658_464# a_534_474# 0.027163f
C26 p2g1 g1 0.007851f
C27 p3 a_594_537# 0.013776f
C28 b1 w_400_n106# 0.015139f
C29 a_594_n65# w_581_n75# 0.019526f
C30 a1 w_548_n81# 0.02809f
C31 w_620_464# g2 0.00583f
C32 a_302_n114# w_328_n116# 0.007992f
C33 c3 w_797_280# 0.012687f
C34 w_238_456# a_218_418# 0.026794f
C35 p1 p1g0 7.17e-19
C36 a_883_464# p3p2g1 3.63e-19
C37 p2 w_538_625# 0.026794f
C38 g2 a_251_466# 0.005106f
C39 p1 a_561_n113# 0.002494f
C40 vdd w_400_28# 0.023245f
C41 a_731_417# a_731_457# 0.41238f
C42 c2 c1 0.013027f
C43 cin g2 0.005207f
C44 vdd a_771_282# 0.019283f
C45 w_604_625# g0 0.026794f
C46 w_642_625# p3p2p1g0 0.013284f
C47 w_660_68# a_597_73# 0.026907f
C48 w_400_28# a_324_88# 0.013216f
C49 w_291_318# a_271_280# 0.026794f
C50 a_825_350# a_883_389# 0.453641f
C51 gnd p2p1g0 0.210726f
C52 w_400_323# a_380_291# 0.026907f
C53 cin w_400_185# 0.00869f
C54 a_873_n248# c2 0.001866f
C55 g2 g1 1.67738f
C56 p0 c3 1.47e-20
C57 w_554_464# a_534_474# 0.027639f
C58 c3 w_867_277# 3.18e-20
C59 vdd a_564_n389# 0.439906f
C60 p2 w_815_n209# 0.028748f
C61 p2 p1 2.60374f
C62 a_561_n113# a1 0.060856f
C63 a_328_n37# a_324_n46# 0.14502f
C64 a_302_n114# a_269_n114# 0.060798f
C65 vdd g3 0.487338f
C66 gnd w_205_450# 2.22e-19
C67 a_738_234# w_725_266# 0.013216f
C68 vdd w_328_n116# 0.001288f
C69 vdd a_518_635# 1.76176f
C70 w_544_301# a_453_311# 0.027163f
C71 p1g0 a_380_291# 0.060798f
C72 w_828_n343# s3 0.015055f
C73 w_400_185# a_380_153# 0.026907f
C74 a_440_393# g0 7.76e-19
C75 w_439_167# a_445_140# 0.008113f
C76 w_439_134# a_445_147# 0.013329f
C77 vdd w_291_180# 6.13e-19
C78 p1 a_534_474# 0.015195f
C79 p2 a_218_418# 0.061185f
C80 cin g0 0.016039f
C81 p0 a_304_190# 0.001371f
C82 p2 w_368_n246# 0.018553f
C83 p3 a_518_635# 0.002444f
C84 cin a_271_142# 0.001372f
C85 p0 pocin 5.46e-21
C86 a_271_142# w_258_174# 0.013216f
C87 c3 w_854_n201# 5.29e-20
C88 gnd a_670_n102# 0.248155f
C89 p3p2p1g0 a_825_350# 0.040556f
C90 vdd a_381_614# 1.32165f
C91 p0 a_302_20# 0.003749f
C92 p1 a_594_n65# 0.004757f
C93 a_594_575# a_518_635# 0.41238f
C94 p2 p3p2p1g0 0.010267f
C95 g1 g0 6.14e-19
C96 p0 p3g2 0.00253f
C97 p1 p3p2g1 0.017215f
C98 a3 g2 0.009821f
C99 p1 a_440_412# 0.013746f
C100 p1 a_610_377# 0.013746f
C101 p3 a_381_614# 0.003255f
C102 pocin a_445_140# 0.185571f
C103 s2 w_854_n201# 0.007992f
C104 vdd a_269_n114# 0.441416f
C105 a_564_n251# vdd 0.439891f
C106 w_347_461# g1 0.01132f
C107 w_725_444# a_731_457# 0.009864f
C108 w_611_272# p1g0 0.001158f
C109 a_798_n113# a_876_n114# 0.14502f
C110 gnd c3 0.42764f
C111 p3 w_368_n380# 0.015055f
C112 vdd b0 0.019072f
C113 a_271_280# g0 0.001372f
C114 a_561_n113# w_548_n81# 0.013216f
C115 a_610_414# a_534_474# 0.41238f
C116 w_584_n351# a_564_n389# 0.026794f
C117 w_660_n346# a_673_n378# 0.013216f
C118 a_594_n65# a1 0.001371f
C119 p1p0c0 a_600_239# 0.211061f
C120 p3g2 p3p2p1p0c0 0.001239f
C121 w_867_n335# p3 0.007896f
C122 p3p2g1 p3p2p1g0 0.0533f
C123 w_328_18# a_302_20# 0.007992f
C124 a_884_498# w_879_518# 0.009864f
C125 a_731_492# w_726_513# 0.009864f
C126 b0 a_324_88# 0.02927f
C127 gnd a_397_472# 0.042086f
C128 a_731_457# a_731_492# 0.41238f
C129 gnd a_304_190# 0.701773f
C130 b3 vdd 0.016782f
C131 b3 w_401_n374# 0.015139f
C132 w_877_451# a_883_429# 0.009864f
C133 g2 w_726_513# 0.036563f
C134 gnd pocin 0.386422f
C135 w_584_n213# b2 0.008451f
C136 p2 a2 0.49284f
C137 w_554_464# p2p1g0 8.56e-21
C138 p1g0 w_400_323# 0.013216f
C139 p0 w_611_340# 1.24e-20
C140 gnd a_302_20# 0.190422f
C141 p3 b3 0.685112f
C142 p1 w_400_n106# 3.76e-36
C143 p1 w_690_n70# 0.002922f
C144 gnd p3g2 0.300358f
C145 p2 a_797_566# 0.013746f
C146 a2 w_329_n250# 0.007896f
C147 p2 c2 0.026943f
C148 gnd a_304_328# 0.588368f
C149 p0 p2g1 0.007444f
C150 p1 p2p1g0 0.016236f
C151 vdd w_551_n357# 0.008823f
C152 b3 a_325_n314# 0.02927f
C153 a_771_282# g3 2.33e-19
C154 p0 w_584_63# 0.00465f
C155 vdd w_879_518# 0.013167f
C156 a_738_234# c2 0.003282f
C157 p2p1p0c0 a_534_474# 0.060798f
C158 a_847_245# w_867_277# 0.026907f
C159 p3 a_797_547# 0.013746f
C160 c2 a_816_233# 3.8e-19
C161 b1 w_367_n112# 0.01395f
C162 a1 w_400_n106# 0.028034f
C163 w_587_464# g2 0.00583f
C164 a_876_n114# c1 0.001856f
C165 a_302_n114# w_291_n117# 0.027261f
C166 a_798_n113# c3 0.001329f
C167 w_205_450# a_218_418# 0.013216f
C168 b3 w_584_n351# 0.008451f
C169 p1 a_670_n102# 0.002494f
C170 a_673_36# w_660_68# 0.013216f
C171 a_564_25# w_584_63# 0.026794f
C172 p0 g2 0.003698f
C173 vdd w_604_625# 0.008451f
C174 vdd a_617_318# 0.41238f
C175 p2 w_521_464# 0.026794f
C176 vdd w_834_277# 0.008512f
C177 cin w_367_185# 0.00869f
C178 p3p2p1p0c0 w_845_654# 0.013216f
C179 p1p0c0 g0 0.010775f
C180 gnd a_600_239# 0.829424f
C181 w_584_63# a_597_73# 0.019526f
C182 w_551_57# a0 0.028093f
C183 w_400_28# b0 0.015139f
C184 w_258_312# a_271_280# 0.013216f
C185 w_367_323# a_380_291# 0.013216f
C186 vdd w_620_464# 0.008451f
C187 gnd p2g1 0.215208f
C188 w_521_464# a_534_474# 0.017642f
C189 vdd a_673_n378# 0.441438f
C190 p2 w_782_n215# 0.028034f
C191 a_380_153# w_367_185# 0.013216f
C192 a_328_n37# b1 0.001802f
C193 a_302_n114# a_324_n46# 0.286223f
C194 a_561_n113# a_594_n65# 0.003752f
C195 s1 w_818_n75# 0.015055f
C196 vdd a_251_466# 0.019451f
C197 gnd a_847_245# 0.248155f
C198 vdd w_291_n117# 0.008507f
C199 vdd a_688_664# 2.20188f
C200 a_251_466# a_327_429# 0.060798f
C201 w_544_301# p1g0 0.004305f
C202 w_506_301# a_453_311# 0.027639f
C203 s2 w_815_n209# 0.015055f
C204 cin vdd 0.057285f
C205 s0 c3 0.003003f
C206 w_611_272# a_617_278# 0.017071f
C207 vdd w_258_174# 0.009216f
C208 w_676_271# a_600_239# 0.027289f
C209 p1 a_397_472# 0.017711f
C210 p2 a_534_474# 0.002444f
C211 p0 g0 0.011127f
C212 w_314_461# a_251_466# 0.026907f
C213 p2 w_329_n250# 0.011491f
C214 p1 w_857_n67# 0.007896f
C215 p3 a_688_664# 0.002444f
C216 p0 a_271_142# 0.060798f
C217 vdd w_807_654# 0.008451f
C218 p3 cin 0.00353f
C219 b3 a_564_n389# 0.00288f
C220 vdd a_380_153# 0.443425f
C221 vdd g1 0.886292f
C222 p3p2g1 a_825_350# 0.001345f
C223 p0 a_269_20# 0.06476f
C224 gnd g2 0.865274f
C225 g1 a_327_429# 0.009049f
C226 p2p1g0 p2p1p0c0 0.057637f
C227 p2 p3p2g1 0.017215f
C228 p1 p3g2 0.057343f
C229 a_738_234# a_816_233# 0.14502f
C230 g0 a_445_140# 0.016231f
C231 a_597_n341# g2 0.013288f
C232 p3p2g1 w_472_604# 0.013216f
C233 c3 c1 2.14e-19
C234 p1 a_304_328# 0.04464f
C235 w_314_461# g1 0.01132f
C236 p2 a_440_412# 0.011867f
C237 p2 a_610_377# 0.013746f
C238 pocin a_445_147# 1.39e-20
C239 p3 g1 0.658617f
C240 p0 w_473_301# 0.026996f
C241 vdd a_324_n46# 0.450999f
C242 w_725_411# p2p1p0c0 0.001174f
C243 vdd w_877_451# 0.010901f
C244 a_798_n113# s1 0.286223f
C245 w_611_305# p1g0 0.036784f
C246 vdd w_367_22# 6.13e-19
C247 vdd a_271_280# 0.455487f
C248 w_942_382# c4 0.013216f
C249 p3 w_329_n384# 0.007992f
C250 gnd a_206_556# 0.20619f
C251 g2 b2 0.764942f
C252 vdd a0 0.236105f
C253 a_873_n248# c3 4.29e-20
C254 w_551_n357# a_564_n389# 0.013216f
C255 p0 a_693_378# 6.43e-21
C256 w_857_n67# c1 0.027735f
C257 p1g0 a_617_278# 0.004158f
C258 a_795_n247# gnd 0.206673f
C259 p3g2 p3p2p1g0 0.001431f
C260 w_828_n343# p3 0.028748f
C261 w_291_17# a_302_20# 0.027261f
C262 g3 w_879_518# 0.036563f
C263 a0 a_324_88# 0.060798f
C264 gnd g0 0.216444f
C265 a_873_n248# s2 0.20619f
C266 b3 w_368_n380# 0.01395f
C267 a3 vdd 0.207557f
C268 a3 w_401_n374# 0.028034f
C269 a_883_429# p3p2p1p0c0 0.005194f
C270 g2 w_658_464# 0.005833f
C271 gnd a_271_142# 0.20619f
C272 w_521_464# p2p1g0 1.11e-19
C273 p1 s1 0.413834f
C274 a_304_328# a_380_291# 0.060798f
C275 w_834_277# a_771_282# 0.027261f
C276 p3 a3 0.413834f
C277 gnd a_269_20# 0.248155f
C278 p1 w_657_n70# 0.002922f
C279 vdd a_325_n180# 0.443244f
C280 c3 c2 0.026004f
C281 w_417_462# g1 2.78e-19
C282 p1 p2g1 0.03968f
C283 p2 p2p1g0 0.001781f
C284 a3 a_325_n314# 0.060798f
C285 w_790_410# c3 0.013216f
C286 s2 c2 0.686118f
C287 w_834_277# g3 0.016049f
C288 p0 w_551_57# 0.00465f
C289 vdd w_726_513# 0.013119f
C290 w_604_625# a_518_635# 0.027639f
C291 a_886_n382# c3 0.002154f
C292 cin a_771_282# 0.68509f
C293 a_693_378# gnd 1.08291f
C294 p2 w_205_450# 0.028034f
C295 p2p1g0 a_534_474# 0.043704f
C296 p3 a_594_556# 0.016756f
C297 a1 w_367_n112# 0.028748f
C298 w_554_464# g2 0.0039f
C299 p3 w_726_513# 4.5e-19
C300 a_673_n378# g3 0.060798f
C301 s1 c1 0.686034f
C302 a_797_566# p3g2 0.004452f
C303 vdd w_708_654# 0.008451f
C304 a_594_556# a_594_575# 0.41238f
C305 s0 a_847_245# 0.060798f
C306 a_597_n341# w_660_n346# 0.026907f
C307 p1 a_328_n37# 6.43e-21
C308 a_564_25# w_551_57# 0.013216f
C309 a_883_429# a_883_464# 0.41238f
C310 a_731_417# p2p1p0c0 0.004158f
C311 a_610_414# p2g1 0.019171f
C312 p1 g2 0.006367f
C313 w_878_485# p3p2p1p0c0 0.018136f
C314 vdd p1p0c0 0.439883f
C315 vdd w_571_625# 0.008451f
C316 vdd w_797_280# 0.001288f
C317 cin w_291_180# 0.008451f
C318 p2 w_401_604# 0.026996f
C319 w_400_28# a0 0.028034f
C320 g3 g1 0.023266f
C321 vdd w_587_464# 0.008451f
C322 c3 a_825_350# 2.29e-19
C323 g2 a_218_418# 0.002036f
C324 a_670_n102# a_594_n65# 0.060798f
C325 a_302_n114# b1 0.685112f
C326 a_594_556# a_594_537# 0.41238f
C327 vdd w_258_n117# 0.008451f
C328 p3p2p1p0c0 a_884_498# 0.005507f
C329 a_269_n114# w_291_n117# 0.013216f
C330 w_506_301# p1g0 0.004305f
C331 w_504_133# g0 0.011197f
C332 w_473_301# a_453_311# 0.027639f
C333 w_795_n349# a_808_n381# 0.013216f
C334 p3 a_329_n305# 0.20619f
C335 s1 c2 0.002762f
C336 w_693_68# g0 0.01325f
C337 p0 vdd 0.810012f
C338 w_611_272# a_600_239# 0.013329f
C339 w_439_134# pocin 1.21e-19
C340 p2 s2 0.413834f
C341 vdd w_867_277# 0.008451f
C342 w_611_305# a_617_278# 0.008113f
C343 a_731_457# w_725_479# 0.009864f
C344 g1 a_381_614# 0.059029f
C345 p1 g0 0.057312f
C346 p3 a_424_535# 0.013746f
C347 p2 a_397_472# 0.002835f
C348 gnd a_808_n381# 0.206673f
C349 vdd w_774_654# 0.008451f
C350 p3 p0 0.002227f
C351 gnd a_302_n114# 0.190422f
C352 p2 w_384_462# 0.026794f
C353 p0 a_324_88# 0.0179f
C354 w_440_301# a_453_311# 0.017642f
C355 a_325_n314# a_329_n305# 0.14502f
C356 a3 a_564_n389# 0.060856f
C357 a_600_239# c2 0.060798f
C358 p3g2 a_825_350# 0.001345f
C359 vdd w_401_n240# 0.026104f
C360 gnd a_239_604# 0.248155f
C361 vdd a_445_140# 0.41238f
C362 p2 p3g2 0.026294f
C363 p2g1 p2p1p0c0 0.008706f
C364 a_883_429# a_883_389# 0.41238f
C365 g0 a_445_147# 0.216537f
C366 cin a_797_585# 2.05e-21
C367 vdd a_564_25# 0.439891f
C368 vdd b1 0.019028f
C369 w_725_444# p2p1p0c0 0.036782f
C370 w_878_485# a_883_464# 0.009864f
C371 vdd p3p2p1p0c0 0.460861f
C372 a_673_36# g0 0.060812f
C373 w_877_383# p3p2p1p0c0 0.053825f
C374 vdd w_328_18# 0.001288f
C375 vdd c4 0.439883f
C376 gnd a_315_567# 0.248155f
C377 w_795_n349# vdd 0.008639f
C378 g2 a2 0.012963f
C379 vdd a_597_73# 0.015633f
C380 a_380_291# g0 0.008577f
C381 a_440_412# a_397_472# 0.41238f
C382 a_670_n102# w_690_n70# 0.026907f
C383 a_239_604# w_302_599# 0.026907f
C384 g2 w_226_594# 0.018971f
C385 p1 w_440_301# 0.026794f
C386 a_302_20# a_328_97# 0.20619f
C387 g0 c1 0.031415f
C388 p1g0 a_600_239# 0.040556f
C389 w_367_22# b0 0.01395f
C390 p3g2 p3p2g1 0.633236f
C391 w_795_n349# p3 0.028034f
C392 vdd gnd 3.52367f
C393 w_291_17# a_269_20# 0.013216f
C394 a0 b0 0.539271f
C395 gnd a_327_429# 0.248155f
C396 a_883_464# a_884_498# 0.41238f
C397 b3 w_329_n384# 0.027716f
C398 a3 w_368_n380# 0.028748f
C399 a_873_n248# a_795_n247# 0.14502f
C400 a_597_n341# vdd 0.011744f
C401 c3 a_876_n114# 6.44e-19
C402 a_883_429# p3p2p1g0 0.00801f
C403 p2p1p0c0 g2 0.065766f
C404 g2 w_193_588# 0.009535f
C405 cin a_797_547# 2.48e-20
C406 w_551_n219# a2 0.028079f
C407 a_206_556# w_226_594# 0.026794f
C408 a_315_567# w_302_599# 0.013216f
C409 p3 gnd 1.77527f
C410 gnd a_324_88# 0.206673f
C411 w_797_280# a_771_282# 0.007992f
C412 a_886_n382# s3 0.20619f
C413 vdd b2 0.003764f
C414 g2 w_238_456# 0.001868f
C415 vdd w_676_271# 0.008511f
C416 a_797_604# a_797_585# 0.41238f
C417 vdd w_302_599# 0.016007f
C418 a_206_556# w_193_588# 0.013216f
C419 a_325_n314# gnd 0.206673f
C420 vdd w_818_n75# 8.63e-20
C421 vdd w_581_n75# 2.04e-19
C422 p2 p2g1 0.004909f
C423 a3 b3 0.535308f
C424 a_795_n247# c2 0.017003f
C425 w_571_625# a_518_635# 0.027639f
C426 vdd w_658_464# 0.008451f
C427 vdd a_883_464# 0.014511f
C428 p0 a_771_282# 0.413834f
C429 p2p1g0 a_397_472# 0.060798f
C430 p1 w_258_312# 0.028034f
C431 p2g1 a_534_474# 9.1e-19
C432 p3 a_424_554# 0.025115f
C433 a_594_n65# w_657_n70# 0.026907f
C434 w_521_464# g2 0.00583f
C435 cin w_620_464# 0.026794f
C436 vdd w_675_654# 0.008451f
C437 w_400_323# g0 0.011443f
C438 a_617_318# g1 0.010567f
C439 a_594_537# gnd 0.412628f
C440 a3 w_551_n357# 0.02808f
C441 a_597_n341# w_584_n351# 0.019526f
C442 p1 a_302_n114# 0.007287f
C443 p3 w_675_654# 0.026794f
C444 cin a_688_664# 0.059029f
C445 p2 g2 0.077377f
C446 w_878_485# p3p2p1g0 0.011197f
C447 vdd w_538_625# 0.008451f
C448 vdd a_453_311# 1.32165f
C449 vdd w_758_272# 6.13e-19
C450 vdd a_798_n113# 0.442386f
C451 p1g0 g0 0.015977f
C452 a_731_417# w_725_411# 0.017071f
C453 w_807_654# a_688_664# 0.027639f
C454 w_367_323# a_304_328# 0.026907f
C455 a_251_466# g1 0.770057f
C456 vdd w_554_464# 0.008451f
C457 cin w_807_654# 0.026794f
C458 s1 a_876_n114# 0.20619f
C459 g2 a_534_474# 0.009442f
C460 a_693_378# p2p1p0c0 0.040556f
C461 cin g1 0.016729f
C462 cin a_380_153# 0.003392f
C463 vdd w_725_266# 0.008698f
C464 a_302_n114# a1 0.413834f
C465 gnd a_771_282# 0.190422f
C466 w_504_133# vdd 0.008451f
C467 a_693_378# w_790_410# 0.027289f
C468 s2 c3 0.015855f
C469 p3p2p1p0c0 g3 0.001229f
C470 vdd w_693_68# 0.008451f
C471 p3p2p1g0 a_884_498# 0.016011f
C472 a_269_n114# w_258_n117# 0.026907f
C473 w_439_134# g0 0.051057f
C474 b1 w_328_n116# 0.027716f
C475 w_473_301# p1g0 0.004305f
C476 w_942_382# a_825_350# 0.027289f
C477 w_877_383# a_883_389# 0.017071f
C478 vdd w_815_n209# 4.8e-19
C479 a_795_n247# w_782_n215# 0.013216f
C480 w_439_167# pocin 0.036563f
C481 p1 vdd 0.796513f
C482 p2 a_795_n247# 0.060798f
C483 w_488_462# p2p1g0 0.013216f
C484 p2 g0 0.033881f
C485 vdd w_505_625# 0.008451f
C486 gnd a_564_n389# 0.20619f
C487 vdd w_741_654# 0.008451f
C488 p3 p1 0.040972f
C489 w_440_301# p1g0 0.004305f
C490 p0 b0 0.023585f
C491 a_597_n341# a_564_n389# 0.003752f
C492 b3 a_329_n305# 0.001802f
C493 vdd a_218_418# 0.439891f
C494 a_600_239# a_617_278# 0.453641f
C495 gnd g3 0.253819f
C496 vdd s0 0.439883f
C497 p3 w_505_625# 0.026794f
C498 gnd a_518_635# 0.042086f
C499 vdd a_445_147# 0.001532f
C500 a_797_604# a_688_664# 0.41238f
C501 p2g1 p2p1g0 0.005273f
C502 p1 a_594_575# 0.031835f
C503 cin a_797_604# 0.013759f
C504 p0 a_797_585# 0.013746f
C505 w_384_462# a_397_472# 0.017642f
C506 vdd a_673_36# 0.441647f
C507 vdd a1 0.230834f
C508 w_725_411# p2g1 0.049155f
C509 vdd p3p2p1g0 0.4601f
C510 w_877_383# p3p2p1g0 0.001142f
C511 w_877_416# p3p2p1p0c0 0.018361f
C512 p3p2g1 g0 0.011924f
C513 vdd w_291_17# 0.008507f
C514 vdd a_380_291# 0.441416f
C515 gnd a_381_614# 0.042086f
C516 p3 p3p2p1g0 0.010267f
C517 w_544_301# g0 0.00229f
C518 vdd c1 0.444335f
C519 a_564_25# b0 0.00288f
C520 a_440_412# g0 0.014522f
C521 a_670_n102# w_657_n70# 0.013216f
C522 a_239_604# w_226_594# 0.019526f
C523 w_328_18# b0 0.027757f
C524 w_367_22# a0 0.028748f
C525 a_564_n251# gnd 0.20619f
C526 gnd a_269_n114# 0.248155f
C527 w_258_17# a_269_20# 0.026907f
C528 a_597_73# b0 0.756776f
C529 p2p1g0 a_731_492# 3.63e-19
C530 a3 w_329_n384# 0.007896f
C531 c3 s1 0.003481f
C532 p2p1g0 g2 0.005084f
C533 p1 w_417_462# 0.026996f
C534 cin w_726_513# 0.002754f
C535 gnd b0 0.045026f
C536 w_758_272# a_771_282# 0.015055f
C537 a_886_n382# a_808_n381# 0.14502f
C538 a_424_554# a_381_614# 0.41238f
C539 a_329_n171# a_325_n180# 0.14502f
C540 a_564_n251# b2 0.002958f
C541 g2 w_205_450# 0.001868f
C542 vdd a2 0.197233f
C543 w_708_654# a_688_664# 0.027639f
C544 vdd w_226_594# 6.13e-19
C545 w_488_462# a_397_472# 0.027163f
C546 s1 w_857_n67# 0.007992f
C547 b3 gnd 0.035921f
C548 vdd w_548_n81# 0.0086f
C549 vdd w_785_n81# 0.030269f
C550 a_597_n341# b3 0.756931f
C551 vdd c2 0.442422f
C552 w_538_625# a_518_635# 0.027639f
C553 c3 a_847_245# 0.006337f
C554 vdd w_193_588# 0.0086f
C555 vdd p2p1p0c0 0.439883f
C556 p3p2p1p0c0 w_879_518# 0.015324f
C557 cin p1p0c0 0.013387f
C558 p2g1 a_397_472# 0.009943f
C559 cin w_797_280# 0.027729f
C560 vdd w_790_410# 0.008495f
C561 p3 w_193_588# 0.028034f
C562 w_384_462# p2g1 1.09e-20
C563 vdd w_400_323# 0.008451f
C564 vdd w_238_456# 6.13e-19
C565 vdd w_642_625# 0.008451f
C566 c3 s3 0.692464f
C567 w_367_323# g0 0.011382f
C568 p1p0c0 g1 0.002848f
C569 a_797_547# gnd 0.41238f
C570 p1 g3 0.028063f
C571 w_584_n213# g2 0.019526f
C572 a_731_417# p2g1 0.019622f
C573 p0 a_688_664# 0.005763f
C574 p1 a_518_635# 0.005763f
C575 vdd p1g0 0.451968f
C576 w_878_485# p3p2g1 6.13e-19
C577 vdd a_561_n113# 0.439891f
C578 p0 cin 0.257529f
C579 p0 w_258_174# 0.028034f
C580 a_518_635# w_505_625# 0.017642f
C581 a_731_417# w_725_444# 0.008113f
C582 w_774_654# a_688_664# 0.027639f
C583 w_291_318# a_304_328# 0.019526f
C584 vdd w_521_464# 0.008451f
C585 g2 a_397_472# 0.00724f
C586 a_693_378# p2p1g0 0.001345f
C587 cin a_496_232# 0.024151f
C588 p0 g1 0.031532f
C589 w_384_462# g2 0.005809f
C590 a_693_378# w_725_411# 0.013329f
C591 vdd a_825_350# 0.011869f
C592 p3p2p1g0 g3 0.001198f
C593 a_795_n247# c3 4.01e-19
C594 a1 w_328_n116# 0.007896f
C595 w_439_167# g0 4.29e-19
C596 vdd w_782_n215# 0.019776f
C597 w_877_383# a_825_350# 0.013329f
C598 w_877_416# a_883_389# 0.008113f
C599 p3p2p1g0 a_518_635# 0.060798f
C600 p3p2p1p0c0 a_688_664# 0.060798f
C601 p1 a_269_n114# 0.06333f
C602 p2 vdd 0.754212f
C603 w_400_185# pocin 0.013216f
C604 g3 c1 0.003696f
C605 vdd w_472_604# 0.008451f
C606 gnd a_673_n378# 0.248155f
C607 a_795_n247# s2 0.286223f
C608 p3 p2 0.395341f
C609 p0 a0 0.007613f
C610 a_597_n341# a_673_n378# 0.060798f
C611 vdd a_534_474# 1.76176f
C612 b1 g1 0.281479f
C613 gnd a_251_466# 0.701773f
C614 vdd a_738_234# 0.439891f
C615 gnd a_440_393# 0.41811f
C616 gnd a_688_664# 0.042086f
C617 g0 a_397_472# 0.059421f
C618 p1 a_797_585# 0.013746f
C619 cin gnd 0.067929f
C620 p0 a_797_604# 0.013746f
C621 a_304_190# a_271_142# 0.003752f
C622 vdd a_594_n65# 0.013824f
C623 a_771_282# c2 0.020436f
C624 vdd p3p2g1 0.454731f
C625 b1 a_324_n46# 0.02927f
C626 w_877_416# p3p2p1g0 0.03763f
C627 w_877_451# p3p2p1p0c0 0.018013f
C628 p3g2 g0 7.61e-19
C629 vdd w_258_17# 0.008451f
C630 vdd w_544_301# 0.008451f
C631 gnd g1 0.512437f
C632 gnd a_380_153# 0.248155f
C633 w_488_462# g2 0.005809f
C634 a_693_378# c3 0.060798f
C635 a_564_25# a0 0.060867f
C636 a_328_97# a_324_88# 0.14502f
C637 a_304_328# g0 0.753587f
C638 p3 p3p2g1 0.017448f
C639 a_269_20# a_302_20# 0.060798f
C640 w_328_18# a0 0.007896f
C641 gnd a_324_n46# 0.206673f
C642 a_594_575# p3p2g1 7.98e-19
C643 g3 c2 0.005387f
C644 a_597_73# a0 0.001371f
C645 p2 a_594_537# 0.020283f
C646 p2g1 g2 0.00516f
C647 cin a_496_251# 0.014005f
C648 gnd a_271_280# 0.20619f
C649 b2 g1 7.83e-19
C650 w_676_271# g1 0.002127f
C651 a_325_n180# w_401_n240# 0.013216f
C652 gnd a0 1.47749f
C653 a_564_n251# a2 0.060856f
C654 a_329_n171# b2 0.001802f
C655 a_424_554# g1 0.013746f
C656 w_675_654# a_688_664# 0.017642f
C657 w_642_625# a_518_635# 0.027163f
C658 w_450_462# a_397_472# 0.027639f
C659 a3 gnd 0.417128f
C660 vdd w_400_n106# 0.026082f
C661 vdd w_690_n70# 0.008451f
C662 a_693_378# a_731_417# 0.453641f
C663 a_597_n341# a3 0.001371f
C664 vdd p2p1g0 0.439883f
C665 w_877_451# a_883_464# 0.01128f
C666 p3p2p1g0 w_879_518# 0.011197f
C667 cin a_453_311# 0.069062f
C668 gnd a_325_n180# 0.206673f
C669 p0 w_797_280# 0.007968f
C670 p2g1 g0 0.002352f
C671 cin w_758_272# 0.013523f
C672 vdd w_660_68# 0.02492f
C673 w_347_461# p2g1 0.013223f
C674 c3 a_808_n381# 0.017003f
C675 vdd w_205_450# 0.0086f
C676 vdd w_367_323# 0.008493f
C677 p0 w_587_464# 0.026996f
C678 a_797_566# a_797_585# 0.41238f
C679 w_291_318# g0 0.008451f
C680 a_738_234# a_771_282# 0.286223f
C681 a_825_350# g3 0.001813f
C682 a_771_282# a_816_233# 0.20619f
C683 p2 g3 0.022389f
C684 b2 a_325_n180# 0.02927f
C685 g2 a_206_556# 0.008991f
C686 p2 a_518_635# 0.004034f
C687 p1 a_440_393# 0.013746f
C688 p0 a_610_395# 0.019134f
C689 p1 a_688_664# 0.004034f
C690 w_878_485# p3g2 0.036563f
C691 vdd a_670_n102# 0.441416f
C692 p1 cin 0.034484f
C693 w_741_654# a_688_664# 0.027639f
C694 a_251_466# a_218_418# 0.003752f
C695 p0 w_774_654# 0.026996f
C696 g2 g0 5.89e-19
C697 a_693_378# p2g1 0.244568f
C698 vdd w_401_604# 0.008451f
C699 p1 g1 0.015873f
C700 a_304_190# w_367_185# 0.026907f
C701 p2 a_381_614# 0.005763f
C702 p0 a_496_232# 0.013746f
C703 w_347_461# g2 0.005799f
C704 w_439_167# vdd 0.0112f
C705 gnd p1p0c0 0.207724f
C706 a_797_566# a_797_547# 0.41238f
C707 w_472_604# a_381_614# 0.027163f
C708 p3g2 a_884_498# 3.63e-19
C709 vdd c3 0.446488f
C710 p3p2g1 g3 0.010274f
C711 p3p2p1g0 a_688_664# 0.00431f
C712 p3p2g1 a_518_635# 0.041586f
C713 p2 a_564_n251# 0.002692f
C714 p0 a_564_25# 0.003966f
C715 p1 a_324_n46# 0.008083f
C716 g1 a_218_418# 0.012164f
C717 p2p1g0 w_725_479# 0.036563f
C718 cin p3p2p1g0 0.02473f
C719 p3g2 w_335_599# 0.013277f
C720 p3 c3 0.03105f
C721 vdd w_434_604# 0.008451f
C722 cin a_610_414# 0.013746f
C723 p1 a_271_280# 0.060798f
C724 p0 a_597_73# 0.007562f
C725 vdd a_397_472# 1.32165f
C726 gnd a_424_535# 0.416913f
C727 a1 g1 0.115698f
C728 vdd a_304_190# 0.017997f
C729 p3g2 a_315_567# 0.060798f
C730 vdd pocin 0.440403f
C731 p3p2g1 a_381_614# 0.060798f
C732 a_693_378# g2 1.39e-20
C733 p0 gnd 0.912787f
C734 vdd w_384_462# 0.008451f
C735 vdd a_302_20# 0.019283f
C736 g1 c1 0.008592f
C737 vdd p3g2 0.447846f
C738 a1 a_324_n46# 0.060798f
C739 w_834_277# c2 8.35e-21
C740 w_877_451# p3p2p1g0 0.012016f
C741 vdd a_304_328# 0.017291f
C742 vdd w_506_301# 0.008451f
C743 gnd a_496_232# 0.41238f
C744 w_450_462# g2 0.005809f
C745 a_302_20# a_324_88# 0.286223f
C746 a_564_25# a_597_73# 0.003752f
C747 a_328_97# b0 0.001802f
C748 p3 p3g2 0.026608f
C749 a_302_n114# w_367_n112# 0.015055f
C750 a_424_554# a_424_535# 0.41238f
C751 gnd a_564_25# 0.20619f
C752 gnd b1 0.03874f
C753 a_797_585# p3p2g1 0.049949f
C754 a_594_575# p3g2 0.042464f
C755 gnd p3p2p1p0c0 0.216485f
C756 a_797_604# p3p2p1g0 0.043431f
C757 p1 a_594_556# 0.018694f
C758 cin a_797_566# 2.14e-20
C759 p2 a_797_547# 0.013746f
C760 gnd c4 0.302435f
C761 a2 g1 0.011016f
C762 p0 a_496_251# 0.013746f
C763 cin c2 0.003312f
C764 b2 w_401_n240# 0.015139f
C765 p1g0 a_617_318# 4.37e-21
C766 a_453_311# p1p0c0 0.060798f
C767 cin p2p1p0c0 0.006726f
C768 gnd a_597_73# 0.248155f
C769 vdd w_693_n346# 0.008611f
C770 a_251_466# w_238_456# 0.019526f
C771 vdd w_488_462# 0.008451f
C772 vdd w_611_340# 0.066855f
C773 w_417_462# a_397_472# 0.027639f
C774 c2 g1 0.014621f
C775 a_496_232# a_496_251# 0.41238f
C776 w_450_462# g0 0.026794f
C777 a_808_n381# s3 0.286223f
C778 a_597_n341# gnd 0.701814f
C779 vdd w_657_n70# 0.008534f
C780 vdd w_367_n112# 6.13e-19
C781 b1 w_581_n75# 0.009938f
C782 a_302_n114# a_328_n37# 0.20619f
C783 c3 a_771_282# 0.007917f
C784 vdd a_600_239# 0.001532f
C785 vdd p2g1 0.439883f
C786 w_238_456# g1 0.021496f
C787 p3p2g1 w_879_518# 4.09e-19
C788 a_883_464# p3p2p1p0c0 0.005542f
C789 p0 a_453_311# 0.005763f
C790 p1 w_571_625# 0.026996f
C791 cin p1g0 0.012177f
C792 p2g1 a_327_429# 0.060798f
C793 gnd b2 0.039673f
C794 p0 w_758_272# 0.028748f
C795 a_239_604# g2 0.75303f
C796 vdd w_584_63# 2.04e-19
C797 vdd w_845_654# 0.008451f
C798 vdd a_847_245# 0.441416f
C799 vdd w_291_318# 6.13e-19
C800 p1g0 g1 0.038781f
C801 c3 g3 0.073145f
C802 p0 w_725_266# 0.028034f
C803 p2 a_251_466# 0.001371f
C804 a2 a_325_n180# 0.060798f
C805 a_239_604# a_206_556# 0.003752f
C806 w_620_464# a_534_474# 0.027639f
C807 p1 w_258_n117# 0.013216f
C808 p1 a_610_395# 0.013746f
C809 p0 w_693_68# 0.001671f
C810 p2 a_440_393# 0.013746f
C811 p2 a_688_664# 0.004034f
C812 p2 cin 0.005346f
C813 w_401_604# a_381_614# 0.027639f
C814 p1 p0 0.069366f
C815 vdd a_731_492# 0.41238f
C816 vdd g2 0.072375f
C817 p3 s3 0.413834f
C818 g2 a_327_429# 0.002808f
C819 vdd w_368_604# 0.008451f
C820 cin a_534_474# 0.060518f
C821 cin a_738_234# 0.024367f
C822 p1 a_496_232# 0.013746f
C823 p2 g1 0.146262f
C824 a_304_190# w_291_180# 0.019526f
C825 s0 w_867_277# 0.013216f
C826 p3 g2 0.017978f
C827 w_314_461# g2 0.005799f
C828 p0 a_445_147# 2.69e-20
C829 w_400_185# vdd 0.02411f
C830 cin a_816_233# 0.002154f
C831 gnd a_453_311# 0.042086f
C832 w_434_604# a_381_614# 0.027639f
C833 gnd a_798_n113# 0.206673f
C834 p3g2 g3 0.013767f
C835 p3 w_368_604# 0.026794f
C836 vdd a_206_556# 0.439891f
C837 vdd w_551_n219# 0.008518f
C838 a_564_n251# w_584_n213# 0.026794f
C839 p3p2p1p0c0 a_883_389# 0.016619f
C840 p3g2 a_518_635# 8.1e-19
C841 p0 a_673_36# 0.003088f
C842 p2 a_329_n171# 0.20619f
C843 w_417_462# p2g1 8.35e-22
C844 p1 b1 0.022716f
C845 cin p3p2g1 0.004802f
C846 p0 p3p2p1g0 0.013325f
C847 p2p1p0c0 a_731_457# 4.37e-21
C848 a_440_412# a_440_393# 0.41238f
C849 a_610_414# a_610_395# 0.41238f
C850 w_867_n335# c3 0.027759f
C851 p3 a_206_556# 0.069923f
C852 vdd a_795_n247# 0.446951f
C853 p0 a_610_414# 0.019134f
C854 a_445_147# a_445_140# 0.453641f
C855 vdd w_942_382# 0.00851f
C856 p0 c1 0.015446f
C857 vdd g0 0.618074f
C858 w_611_272# p1p0c0 0.057514f
C859 w_611_305# a_617_318# 0.009864f
C860 p3g2 a_381_614# 0.011947f
C861 vdd a_271_142# 0.439904f
C862 vdd w_347_461# 0.008451f
C863 p1 gnd 0.59676f
C864 w_347_461# a_327_429# 0.026907f
C865 vdd a_269_20# 0.441416f
C866 a1 b1 0.614689f
C867 a_617_318# a_617_278# 0.41238f
C868 a_453_311# a_496_251# 0.41238f
C869 w_693_n346# g3 0.013222f
C870 w_877_451# p3p2g1 0.037044f
C871 p3p2p1g0 p3p2p1p0c0 0.003212f
C872 w_797_280# c2 0.003455f
C873 gnd a_218_418# 0.208267f
C874 vdd w_473_301# 0.008451f
C875 vdd a_883_429# 5.02e-19
C876 a_594_575# g0 0.013746f
C877 a_731_492# w_725_479# 0.01128f
C878 gnd s0 0.20619f
C879 w_417_462# g2 0.005809f
C880 a_673_36# a_597_73# 0.060798f
C881 a_302_20# b0 0.685117f
C882 gnd a_445_147# 0.576829f
C883 w_620_464# p2p1g0 9.19e-21
C884 p2 a_325_n180# 0.288532f
C885 a_771_282# a_847_245# 0.060798f
C886 gnd a_673_36# 0.248155f
C887 gnd a1 1.83674f
C888 p1 w_818_n75# 0.028748f
C889 p1 w_581_n75# 0.002922f
C890 vdd w_440_301# 0.008451f
C891 a_797_585# p3g2 0.054573f
C892 gnd p3p2p1g0 0.232346f
C893 a_797_604# p3p2g1 0.003102f
C894 vdd a_693_378# 0.001532f
C895 c1 a_597_73# 2.15e-19
C896 p2 a_594_556# 0.023173f
C897 gnd a_380_291# 0.248155f
C898 p0 c2 0.020959f
C899 b2 w_368_n246# 0.01395f
C900 w_611_305# g1 0.002086f
C901 a2 w_401_n240# 0.028034f
C902 p1g0 p1p0c0 0.011688f
C903 gnd c1 0.261394f
C904 cin p2p1g0 0.070233f
C905 p0 p2p1p0c0 0.00185f
C906 w_878_485# a_884_498# 0.01128f
C907 g1 w_690_n70# 0.01323f
C908 vdd w_660_n346# 0.008611f
C909 g3 a_847_245# 0.015251f
C910 vdd w_450_462# 0.008451f
C911 p2 w_708_654# 0.026794f
C912 a_324_n46# w_400_n106# 0.013216f
C913 c2 w_854_n201# 0.027735f
C914 a_797_547# p3g2 0.001272f
C915 c3 w_834_277# 3.18e-20
C916 w_205_450# g1 0.013044f
C917 w_818_n75# c1 0.015306f
C918 g2 g3 0.005441f
C919 p1 a_453_311# 0.002444f
C920 p0 p1g0 7.17e-19
C921 a_883_464# p3p2p1g0 0.016011f
C922 p1 a_798_n113# 0.060798f
C923 gnd a2 1.55938f
C924 vdd w_551_57# 0.0086f
C925 p1 w_554_464# 0.041309f
C926 vdd w_258_312# 0.028134f
C927 gnd c2 0.219293f
C928 a_670_n102# g1 0.060798f
C929 w_584_63# b0 0.008938f
C930 gnd p2p1p0c0 0.207724f
C931 p2 a_424_535# 0.023137f
C932 a_239_604# a_315_567# 0.060798f
C933 a2 b2 0.531092f
C934 w_587_464# a_534_474# 0.027639f
C935 cin c3 5.08e-19
C936 vdd a_808_n381# 0.439903f
C937 w_368_604# a_381_614# 0.017642f
C938 w_335_599# a_315_567# 0.026907f
C939 vdd a_302_n114# 0.019283f
C940 p2 p0 0.021197f
C941 a_561_n113# b1 0.00343f
C942 vdd a_884_498# 0.41238f
C943 gnd w_238_456# 0.003687f
C944 vdd a_239_604# 0.024911f
C945 a_564_n251# g2 0.003752f
C946 w_544_301# p1p0c0 0.013229f
C947 g3 g0 0.00202f
C948 w_867_n335# s3 0.007992f
C949 p3 a_808_n381# 0.060798f
C950 p1 w_741_654# 0.026794f
C951 a_518_635# g0 0.059018f
C952 vdd w_367_185# 0.008465f
C953 w_504_133# a_445_147# 0.027289f
C954 w_439_134# a_445_140# 0.017071f
C955 w_676_271# c2 0.016933f
C956 vdd w_335_599# 0.008451f
C957 a_798_n113# c1 0.016996f
C958 p0 a_534_474# 0.005763f
C959 p0 a_738_234# 0.060798f
C960 cin a_304_190# 0.747651f
C961 c2 w_818_n75# 0.019549f
C962 p2 w_401_n240# 0.003504f
C963 p3 a_239_604# 0.002112f
C964 cin pocin 0.002387f
C965 a_271_142# w_291_180# 0.026794f
C966 gnd p1g0 0.207724f
C967 w_693_68# a_673_36# 0.026907f
C968 w_434_604# g1 0.026794f
C969 gnd a_561_n113# 0.20619f
C970 p3p2p1p0c0 a_825_350# 0.217915f
C971 p3p2p1g0 a_883_389# 0.004158f
C972 a_564_n251# w_551_n219# 0.013216f
C973 vdd a_315_567# 0.464809f
C974 p0 a_328_97# 3.98e-19
C975 p2 w_854_n201# 0.007896f
C976 p1 a1 0.008941f
C977 p0 p3p2g1 0.012004f
C978 g1 a_397_472# 0.007928f
C979 cin p3g2 0.004802f
C980 p2p1p0c0 w_658_464# 0.013216f
C981 p1 p3p2p1g0 0.010267f
C982 a_304_190# a_380_153# 0.060798f
C983 a_825_350# c4 0.060798f
C984 a_610_395# a_610_377# 0.41238f
C985 b3 g2 3.99e-19
C986 w_504_133# c1 0.013242f
C987 a_380_153# pocin 0.060798f
C988 w_828_n343# c3 0.016729f
C989 p0 w_258_17# 0.013216f
C990 p3 a_315_567# 0.001362f
C991 p0 a_610_377# 6.84e-20
C992 cin w_506_301# 0.026794f
C993 w_384_462# g1 0.011399f
C994 vdd w_401_n374# 0.028764f
C995 p1 c1 0.024407f
C996 vdd a_327_429# 0.441435f
C997 w_611_340# a_617_318# 0.009864f
C998 w_611_305# p1p0c0 1.04e-20
C999 p3g2 g1 0.023512f
C1000 gnd a_825_350# 1.36074f
C1001 vdd w_314_461# 0.012946f
C1002 p3 vdd 0.984731f
C1003 p2 gnd 1.81974f
C1004 vdd a_324_88# 0.45515f
C1005 a_561_n113# w_581_n75# 0.026794f
C1006 a_798_n113# w_785_n81# 0.013216f
C1007 w_693_n346# a_673_n378# 0.026907f
C1008 w_314_461# a_327_429# 0.013216f
C1009 a_594_n65# b1 0.7623f
C1010 p1p0c0 a_617_278# 0.019123f
C1011 w_758_272# c2 0.003448f
C1012 p3p2g1 p3p2p1p0c0 0.001238f
C1013 c1 a_445_147# 0.060798f
C1014 a_798_n113# c2 0.003242f
C1015 w_367_22# a_302_20# 0.015055f
C1016 gnd a_534_474# 0.042086f
C1017 a_325_n314# vdd 0.442574f
C1018 gnd a_738_234# 0.206673f
C1019 a_325_n314# w_401_n374# 0.013216f
C1020 w_877_416# a_883_429# 0.009864f
C1021 a_302_20# a0 0.413834f
C1022 p3 a_594_575# 2.95e-20
C1023 w_587_464# p2p1g0 8.56e-21
C1024 p2 b2 0.6987f
C1025 a_886_n382# 0 0.016528f **FLOATING
C1026 s3 0 0.473154f **FLOATING
C1027 a_808_n381# 0 0.526842f **FLOATING
C1028 a_564_n389# 0 0.477455f **FLOATING
C1029 a_673_n378# 0 0.382299f **FLOATING
C1030 a_329_n305# 0 0.016528f **FLOATING
C1031 a_325_n314# 0 0.526842f **FLOATING
C1032 b3 0 6.62907f **FLOATING
C1033 a3 0 2.45012f **FLOATING
C1034 a_597_n341# 0 0.771781f **FLOATING
C1035 a_873_n248# 0 0.016528f **FLOATING
C1036 s2 0 0.462937f **FLOATING
C1037 a_795_n247# 0 0.526842f **FLOATING
C1038 vdd 0 37.96201f **FLOATING
C1039 a_564_n251# 0 0.477455f **FLOATING
C1040 a_329_n171# 0 0.016528f **FLOATING
C1041 a_325_n180# 0 0.526842f **FLOATING
C1042 b2 0 6.55321f **FLOATING
C1043 a2 0 2.34823f **FLOATING
C1044 a_876_n114# 0 0.016528f **FLOATING
C1045 s1 0 0.462937f **FLOATING
C1046 a_798_n113# 0 0.526842f **FLOATING
C1047 a_561_n113# 0 0.477455f **FLOATING
C1048 a_670_n102# 0 0.382299f **FLOATING
C1049 a_328_n37# 0 0.016528f **FLOATING
C1050 a_302_n114# 0 0.662497f **FLOATING
C1051 a_269_n114# 0 0.382299f **FLOATING
C1052 a_324_n46# 0 0.526842f **FLOATING
C1053 b1 0 5.67351f **FLOATING
C1054 a1 0 2.3497f **FLOATING
C1055 a_594_n65# 0 0.771781f **FLOATING
C1056 a_564_25# 0 0.477455f **FLOATING
C1057 a_673_36# 0 0.382299f **FLOATING
C1058 a_328_97# 0 0.016528f **FLOATING
C1059 a_302_20# 0 0.662497f **FLOATING
C1060 a_269_20# 0 0.382299f **FLOATING
C1061 a_324_88# 0 0.526842f **FLOATING
C1062 b0 0 6.55052f **FLOATING
C1063 a0 0 2.47333f **FLOATING
C1064 a_597_73# 0 0.804448f **FLOATING
C1065 c1 0 2.23371f **FLOATING
C1066 a_445_140# 0 0.179875f **FLOATING
C1067 a_445_147# 0 1.02677f **FLOATING
C1068 a_816_233# 0 0.016528f **FLOATING
C1069 pocin 0 0.599293f **FLOATING
C1070 a_271_142# 0 0.477455f **FLOATING
C1071 a_380_153# 0 0.382299f **FLOATING
C1072 a_496_232# 0 0.040245f **FLOATING
C1073 s0 0 0.145867f **FLOATING
C1074 a_738_234# 0 0.526842f **FLOATING
C1075 a_304_190# 0 0.771781f **FLOATING
C1076 a_496_251# 0 0.040245f **FLOATING
C1077 c2 0 2.27948f **FLOATING
C1078 a_617_278# 0 0.206277f **FLOATING
C1079 a_600_239# 0 1.28245f **FLOATING
C1080 a_847_245# 0 0.382299f **FLOATING
C1081 a_771_282# 0 0.662497f **FLOATING
C1082 a_617_318# 0 0.150155f **FLOATING
C1083 p1p0c0 0 0.596493f **FLOATING
C1084 a_453_311# 0 1.70512f **FLOATING
C1085 p1g0 0 1.48359f **FLOATING
C1086 a_271_280# 0 0.477455f **FLOATING
C1087 c4 0 0.147767f **FLOATING
C1088 a_380_291# 0 0.382299f **FLOATING
C1089 a_610_377# 0 0.036687f **FLOATING
C1090 a_304_328# 0 0.771914f **FLOATING
C1091 a_440_393# 0 0.040245f **FLOATING
C1092 a_610_395# 0 0.040245f **FLOATING
C1093 a_883_389# 0 0.206277f **FLOATING
C1094 a_825_350# 0 1.81542f **FLOATING
C1095 c3 0 2.59712f **FLOATING
C1096 a_610_414# 0 0.040245f **FLOATING
C1097 a_440_412# 0 0.040245f **FLOATING
C1098 a_731_417# 0 0.206277f **FLOATING
C1099 a_883_429# 0 0.150155f **FLOATING
C1100 a_693_378# 0 1.54889f **FLOATING
C1101 a_731_457# 0 0.150155f **FLOATING
C1102 a_883_464# 0 0.148414f **FLOATING
C1103 p2p1p0c0 0 1.73078f **FLOATING
C1104 p2p1g0 0 1.59696f **FLOATING
C1105 p2g1 0 0.842448f **FLOATING
C1106 a_218_418# 0 0.477455f **FLOATING
C1107 a_534_474# 0 2.13082f **FLOATING
C1108 a_397_472# 0 1.70506f **FLOATING
C1109 g0 0 11.784104f **FLOATING
C1110 a_327_429# 0 0.382299f **FLOATING
C1111 a_731_492# 0 0.148414f **FLOATING
C1112 a_884_498# 0 0.144831f **FLOATING
C1113 g3 0 6.00295f **FLOATING
C1114 a_251_466# 0 0.770807f **FLOATING
C1115 a_424_535# 0 0.040245f **FLOATING
C1116 a_594_537# 0 0.040245f **FLOATING
C1117 a_797_547# 0 0.040245f **FLOATING
C1118 a_594_556# 0 0.040245f **FLOATING
C1119 a_424_554# 0 0.040245f **FLOATING
C1120 a_797_566# 0 0.040245f **FLOATING
C1121 a_594_575# 0 0.040245f **FLOATING
C1122 a_797_585# 0 0.040245f **FLOATING
C1123 a_797_604# 0 0.040245f **FLOATING
C1124 gnd 0 32.5503f **FLOATING
C1125 p3p2p1p0c0 0 4.09846f **FLOATING
C1126 p3p2p1g0 0 6.27811f **FLOATING
C1127 p3p2g1 0 4.70971f **FLOATING
C1128 p3g2 0 5.74969f **FLOATING
C1129 a_206_556# 0 0.477455f **FLOATING
C1130 a_315_567# 0 0.382299f **FLOATING
C1131 a_381_614# 0 1.70511f **FLOATING
C1132 g1 0 21.4853f **FLOATING
C1133 g2 0 19.795301f **FLOATING
C1134 a_239_604# 0 0.804448f **FLOATING
C1135 a_518_635# 0 2.1423f **FLOATING
C1136 a_688_664# 0 2.57948f **FLOATING
C1137 cin 0 4.54341f **FLOATING
C1138 p0 0 7.2243f **FLOATING
C1139 p1 0 13.8549f **FLOATING
C1140 p2 0 13.4502f **FLOATING
C1141 p3 0 15.000999f **FLOATING
C1142 w_867_n335# 0 1.25349f **FLOATING
C1143 w_828_n343# 0 1.34991f **FLOATING
C1144 w_795_n349# 0 1.34991f **FLOATING
C1145 w_693_n346# 0 1.34991f **FLOATING
C1146 w_660_n346# 0 1.34991f **FLOATING
C1147 w_584_n351# 0 1.34991f **FLOATING
C1148 w_551_n357# 0 1.34991f **FLOATING
C1149 w_401_n374# 0 1.34991f **FLOATING
C1150 w_368_n380# 0 1.34991f **FLOATING
C1151 w_329_n384# 0 1.25349f **FLOATING
C1152 w_854_n201# 0 1.25349f **FLOATING
C1153 w_815_n209# 0 1.34991f **FLOATING
C1154 w_782_n215# 0 1.34991f **FLOATING
C1155 w_584_n213# 0 1.34991f **FLOATING
C1156 w_551_n219# 0 1.34991f **FLOATING
C1157 w_401_n240# 0 1.34991f **FLOATING
C1158 w_368_n246# 0 1.34991f **FLOATING
C1159 w_329_n250# 0 1.25349f **FLOATING
C1160 w_857_n67# 0 1.25349f **FLOATING
C1161 w_818_n75# 0 1.34991f **FLOATING
C1162 w_785_n81# 0 1.34991f **FLOATING
C1163 w_690_n70# 0 1.34991f **FLOATING
C1164 w_657_n70# 0 1.34991f **FLOATING
C1165 w_581_n75# 0 1.34991f **FLOATING
C1166 w_548_n81# 0 1.34991f **FLOATING
C1167 w_400_n106# 0 1.34991f **FLOATING
C1168 w_367_n112# 0 1.34991f **FLOATING
C1169 w_328_n116# 0 1.25349f **FLOATING
C1170 w_291_n117# 0 1.34991f **FLOATING
C1171 w_258_n117# 0 1.34991f **FLOATING
C1172 w_693_68# 0 1.34991f **FLOATING
C1173 w_660_68# 0 1.34991f **FLOATING
C1174 w_584_63# 0 1.34991f **FLOATING
C1175 w_551_57# 0 1.34991f **FLOATING
C1176 w_400_28# 0 1.34991f **FLOATING
C1177 w_367_22# 0 1.34991f **FLOATING
C1178 w_328_18# 0 1.25349f **FLOATING
C1179 w_291_17# 0 1.34991f **FLOATING
C1180 w_258_17# 0 1.34991f **FLOATING
C1181 w_504_133# 0 1.34991f **FLOATING
C1182 w_439_134# 0 1.34991f **FLOATING
C1183 w_439_167# 0 1.34991f **FLOATING
C1184 w_400_185# 0 1.34991f **FLOATING
C1185 w_367_185# 0 1.34991f **FLOATING
C1186 w_291_180# 0 1.34991f **FLOATING
C1187 w_258_174# 0 1.34991f **FLOATING
C1188 w_867_277# 0 1.34991f **FLOATING
C1189 w_834_277# 0 1.34991f **FLOATING
C1190 w_797_280# 0 1.25349f **FLOATING
C1191 w_758_272# 0 1.34991f **FLOATING
C1192 w_725_266# 0 1.34991f **FLOATING
C1193 w_676_271# 0 1.34991f **FLOATING
C1194 w_611_272# 0 1.34991f **FLOATING
C1195 w_611_305# 0 1.34991f **FLOATING
C1196 w_611_340# 0 1.34991f **FLOATING
C1197 w_544_301# 0 1.34991f **FLOATING
C1198 w_506_301# 0 1.34991f **FLOATING
C1199 w_473_301# 0 1.34991f **FLOATING
C1200 w_440_301# 0 1.34991f **FLOATING
C1201 w_400_323# 0 1.34991f **FLOATING
C1202 w_367_323# 0 1.34991f **FLOATING
C1203 w_291_318# 0 1.34991f **FLOATING
C1204 w_258_312# 0 1.34991f **FLOATING
C1205 w_942_382# 0 1.34991f **FLOATING
C1206 w_877_383# 0 1.34991f **FLOATING
C1207 w_877_416# 0 1.34991f **FLOATING
C1208 w_877_451# 0 1.34991f **FLOATING
C1209 w_790_410# 0 1.34991f **FLOATING
C1210 w_725_411# 0 1.34991f **FLOATING
C1211 w_725_444# 0 1.34991f **FLOATING
C1212 w_878_485# 0 1.34991f **FLOATING
C1213 w_725_479# 0 1.34991f **FLOATING
C1214 w_879_518# 0 1.34991f **FLOATING
C1215 w_726_513# 0 1.34991f **FLOATING
C1216 w_658_464# 0 1.34991f **FLOATING
C1217 w_620_464# 0 1.34991f **FLOATING
C1218 w_587_464# 0 1.34991f **FLOATING
C1219 w_554_464# 0 1.34991f **FLOATING
C1220 w_521_464# 0 1.34991f **FLOATING
C1221 w_488_462# 0 1.34991f **FLOATING
C1222 w_450_462# 0 1.34991f **FLOATING
C1223 w_417_462# 0 1.34991f **FLOATING
C1224 w_384_462# 0 1.34991f **FLOATING
C1225 w_347_461# 0 1.34991f **FLOATING
C1226 w_314_461# 0 1.34991f **FLOATING
C1227 w_238_456# 0 1.34991f **FLOATING
C1228 w_205_450# 0 1.34991f **FLOATING
C1229 w_845_654# 0 1.34991f **FLOATING
C1230 w_807_654# 0 1.34991f **FLOATING
C1231 w_774_654# 0 1.34991f **FLOATING
C1232 w_741_654# 0 1.34991f **FLOATING
C1233 w_708_654# 0 1.34991f **FLOATING
C1234 w_675_654# 0 1.34991f **FLOATING
C1235 w_642_625# 0 1.34991f **FLOATING
C1236 w_604_625# 0 1.34991f **FLOATING
C1237 w_571_625# 0 1.34991f **FLOATING
C1238 w_538_625# 0 1.34991f **FLOATING
C1239 w_505_625# 0 1.34991f **FLOATING
C1240 w_472_604# 0 1.34991f **FLOATING
C1241 w_434_604# 0 1.34991f **FLOATING
C1242 w_401_604# 0 1.34991f **FLOATING
C1243 w_368_604# 0 1.34991f **FLOATING
C1244 w_335_599# 0 1.34991f **FLOATING
C1245 w_302_599# 0 1.34991f **FLOATING
C1246 w_226_594# 0 1.34991f **FLOATING
C1247 w_193_588# 0 1.34991f **FLOATING
