* SPICE3 file created from cla.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Power Supply for the circuit
Vdd vdd gnd 'SUPPLY'


* Input Signals
* for testing
* Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
* Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 30n 60n)     
* Va1 a1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 10n 20n)    
* Vb1 b1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 30n 60n)    
* Va2 a2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 10n 20n)   
* Vb2 b2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 30n 60n)   
* Va3 a3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 10n 20n)   
* Vb3 b3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 30n 60n)   
* Vcin cin gnd DC 0         

* Input Signals for delay measurement
*  rising
Vclk clk gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)  
Va0 a0 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)     
Vb0 b0 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)     
Va1 a1 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)    
Vb1 b1 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)    
Va2 a2 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Vb2 b2 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Va3 a3 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Vb3 b3 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Vcin cin gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)


* Input Signals for delay measurement
*  falling
* Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
* Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Va1 a1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
* Vb1 b1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
* Va2 a2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Vb2 b2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Va3 a3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Vb3 b3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Vcin cin gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)                             





.option scale=0.09u

M1000 a_445_147# g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 a_691_n240# a_615_n203# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_615_n203# a_582_n251# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 p2g1 a_327_429# vdd w_347_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_610_376# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1005 a_594_575# p1 a_594_556# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 a_440_412# p1 a_440_393# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 p1p0c0 a_453_311# vdd w_544_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 a3 a_338_n335# a_303_n382# w_329_n384# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1009 a_848_2# p2 c2 w_835_n8# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_518_635# p3 vdd w_505_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1011 a_731_457# p2p1p0c0 a_731_417# w_725_444# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1012 b2 a2 a_303_n248# w_368_n246# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1013 gnd a_303_n248# a_270_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 p3p2g1 a_381_614# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1015 p2p1p0c0 a_534_474# vdd w_658_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1016 a_610_395# p1 a_610_376# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1017 gnd a_325_n180# a_303_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1018 a_815_n46# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1019 a_518_635# g0 a_594_575# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1020 a_940_n169# a_864_n132# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1021 s2 a_924_n35# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1022 vdd a0 a_345_92# w_400_28# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 vdd a_302_20# a_269_20# w_291_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1024 a_346_n176# b2 a_303_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1025 g0 a_691_36# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1026 a_825_350# p3p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 a_847_245# a_771_282# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1028 a_304_190# a_271_142# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1029 a_884_498# p3g2 a_883_464# w_878_485# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1030 g3 a_691_n378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1031 a_731_492# p2g1g0 a_731_457# w_725_479# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1032 a_831_148# a_879_123# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1033 a_615_n341# a3 b3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1034 a_831_148# a_866_144# p1 w_857_147# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1035 a_798_100# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 a_315_567# a_239_604# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1037 g2 a_691_n240# vdd w_711_n208# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1038 a_582_n251# a2 vdd w_569_n219# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1039 p3g2 a_315_567# vdd w_335_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 vdd g3 a_884_498# w_879_518# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1041 a_825_350# p3p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1042 pocin a_380_153# vdd w_400_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1043 vdd a_269_20# p0 w_258_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1044 a_218_418# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1045 a_380_153# a_304_190# vdd w_367_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 b1 a1 a_302_n114# w_367_n112# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1047 a_691_36# a_615_73# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 a_825_350# p3p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1049 a_271_280# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1050 a_907_111# a_831_148# vdd w_894_143# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1051 s2 a_924_n35# vdd w_944_n3# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 p3p2p1g0 a_518_635# vdd w_642_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_615_n203# a_582_n251# b2 w_602_n213# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1054 a_239_604# a_206_556# g2 w_226_594# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1055 a_304_190# a_271_142# cin w_291_180# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_612_n65# a_579_n113# b1 w_599_n75# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 a_582_25# a0 vdd w_569_57# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 p2p1g0 a_397_472# vdd w_488_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1059 c3 a_693_378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1060 a_440_393# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1061 a_612_n65# a_579_n113# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1062 a_924_n35# a_848_2# vdd w_911_n3# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 a_688_664# p0 vdd w_774_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1064 a_445_147# pocin gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 p2g1 a_327_429# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 a_600_239# p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1067 s3 a_940_n169# vdd w_960_n137# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_327_429# a_251_466# vdd w_314_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1069 a_848_2# a_896_n23# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1070 a_688_664# cin vdd w_807_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1071 a_693_378# p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_251_466# p2 g1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 a_346_n310# b3 a_303_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_688_n102# a_612_n65# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1075 a_738_234# p0 vdd w_725_266# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1076 a_924_n35# a_848_2# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1077 p3p2g1 a_381_614# vdd w_472_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1078 a_206_556# p3 vdd w_193_588# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1079 a_424_535# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1080 g2 a_691_n240# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1081 s0 a_847_245# vdd w_867_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_582_n389# a3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1083 a_691_n378# a_615_n341# vdd w_678_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1084 a_864_n132# a_912_n157# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1085 vdd a2 a_346_n176# w_401_n240# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_615_n203# a2 b2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1087 g1 a_688_n102# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1088 c4 a_825_350# vdd w_942_382# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_424_554# p2 a_424_535# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 a_453_311# p0 vdd w_473_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_831_n180# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_315_567# a_239_604# vdd w_302_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 p3p2p1p0c0 a_688_664# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1094 a_771_282# p0 cin w_758_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 a_271_142# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_612_n65# a1 b1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1097 a_534_474# cin vdd w_620_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_534_474# p0 vdd w_587_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1099 a_453_311# cin vdd w_506_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_271_280# p1 vdd w_258_312# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_693_378# p2g1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1102 a_381_614# g1 a_424_554# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_883_429# p3p2p1g0 a_883_389# w_877_416# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 c1 a_445_147# vdd w_504_133# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_304_328# a_271_280# g0 w_291_318# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_825_350# p3g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 a_688_664# p1 vdd w_741_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_797_604# p0 a_797_585# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 vdd a_269_n114# p1 w_258_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1110 p1g0 a_380_291# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 a_345_n42# b1 a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_327_429# a_251_466# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1113 a1 a_337_n67# a_302_n114# w_328_n116# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 s1 a_907_111# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1115 a_693_378# p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_380_291# a_304_328# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 c2 a_600_239# vdd w_676_271# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1118 gnd a_324_88# a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 b3 a3 a_303_n382# w_368_n380# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1120 a_688_n102# a_612_n65# vdd w_675_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 gnd a_324_n46# a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1122 a_815_n46# p2 vdd w_802_n14# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 vdd a3 a_346_n310# w_401_n374# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1124 a_615_73# a_582_25# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 p1p0c0 a_453_311# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1126 a_345_92# b0 a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 a_688_664# cin a_797_604# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1128 vdd g2 a_731_492# w_726_513# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1129 a_883_464# p3p2g1 a_883_429# w_877_451# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 a_693_378# g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1131 g1 a_688_n102# vdd w_708_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_831_148# c1 a_798_100# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_864_n132# p3 c3 w_851_n142# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1134 a_304_328# p1 g0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1135 a_771_282# a_819_257# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1136 a_518_635# p1 vdd w_571_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1137 a_397_472# g0 vdd w_450_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1138 a_579_n113# a1 vdd w_566_n81# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_797_547# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_496_251# p0 a_496_232# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_848_2# a_883_n2# p2 w_874_1# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 g0 a_691_36# vdd w_711_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_847_245# a_771_282# vdd w_834_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1147 vdd a_270_n248# p2 w_259_n251# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1148 a_579_n113# a1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1149 a_239_604# a_206_556# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1150 a_797_566# p2 a_797_547# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 a_453_311# cin a_496_251# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1152 a_453_311# p1 vdd w_440_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_798_100# p1 vdd w_785_132# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1154 gnd a3 a_346_n310# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1155 a_534_474# p1 vdd w_554_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 a_304_328# a_271_280# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_445_147# g0 a_445_140# w_439_134# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1158 a_940_n169# a_864_n132# vdd w_927_n137# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1159 a_797_585# p1 a_797_566# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1160 a_864_n132# c3 a_831_n180# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1161 gnd a_302_n114# a_269_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_691_36# a_615_73# vdd w_678_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1163 s3 a_940_n169# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_864_n132# a_899_n136# p3 w_890_n133# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1165 gnd a_269_n114# p1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1166 a_381_614# g1 vdd w_434_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1167 vdd a_303_n248# a_270_n248# w_292_n251# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 pocin a_380_153# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 a_848_2# c2 a_815_n46# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1170 a_380_153# a_304_190# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 a_831_148# p1 c1 w_818_138# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1172 a_688_664# p3 vdd w_675_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 g3 a_691_n378# vdd w_711_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_907_111# a_831_148# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1175 p1g0 a_380_291# vdd w_400_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1176 c2 a_600_239# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 a_615_73# a0 b0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1178 a0 a_337_67# a_302_20# w_328_18# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_380_291# a_304_328# vdd w_367_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1180 vdd a_270_n382# p3 w_259_n385# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1181 a_582_25# a0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1182 a_688_664# p2 vdd w_708_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 p2p1g0 a_397_472# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1184 gnd a2 a_346_n176# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1185 vdd pocin a_445_140# w_439_167# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 c3 a_693_378# vdd w_790_410# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1187 a_304_190# p0 cin Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_251_466# a_218_418# g1 w_238_456# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 vdd a1 a_345_n42# w_400_n106# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# g0 a_440_412# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 a_691_n378# a_615_n341# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1192 a_615_n341# a_582_n389# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1193 a_397_472# p2 vdd w_384_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 vdd a_303_n382# a_270_n382# w_292_n385# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1195 vdd a_302_n114# a_269_n114# w_291_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_617_318# p1g0 a_617_278# w_611_305# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 a_771_282# a_806_278# p0 w_797_281# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_738_234# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1199 a_691_n240# a_615_n203# vdd w_678_n208# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_518_635# p2 vdd w_538_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1201 a_496_232# p1 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 b0 a0 a_302_20# w_367_22# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_397_472# p1 vdd w_417_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_206_556# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1205 gnd a_270_n382# p3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 a_610_414# p0 a_610_395# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 p3p2p1p0c0 a_688_664# vdd w_845_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1208 a_271_142# p0 vdd w_258_174# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1209 a_582_n251# a2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 a_534_474# p2 vdd w_521_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1211 s0 a_847_245# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1212 vdd g1 a_617_318# w_611_340# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 c4 a_825_350# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 gnd a0 a_345_92# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1215 gnd a1 a_345_n42# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 gnd a_302_20# a_269_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1217 a_381_614# p2 vdd w_401_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1218 a_534_474# cin a_610_414# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1219 a2 a_338_n201# a_303_n248# w_329_n250# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1220 a_251_466# a_218_418# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1221 a_771_282# cin a_738_234# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1222 a_381_614# p3 vdd w_368_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1223 p3g2 a_315_567# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1224 a_594_537# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1225 a_600_239# g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1226 a_615_73# a_582_25# b0 w_602_63# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1227 a_582_n389# a3 vdd w_569_n357# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1228 a_239_604# p3 g2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1229 gnd a_325_n314# a_303_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1230 gnd a_303_n382# a_270_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1231 a_218_418# p2 vdd w_205_450# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1232 a_825_350# g3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1233 a_600_239# p1p0c0 a_617_278# w_611_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1234 s1 a_907_111# vdd w_927_143# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1235 c1 a_445_147# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1236 p3p2p1g0 a_518_635# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1237 a_693_378# p2g1 a_731_417# w_725_411# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1238 a_831_n180# p3 vdd w_818_n148# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1239 a_600_239# p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1240 gnd a_270_n248# p2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1241 a_594_556# p2 a_594_537# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1242 gnd a_269_20# p0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1243 a_615_n341# a_582_n389# b3 w_602_n351# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 w_877_416# a_883_389# 1.128f
C1 w_942_382# a_825_350# 1.014f
C2 w_329_n250# a_303_n248# 1.128f
C3 w_927_143# s1 1.88f
C4 w_774_654# p0 1.014f
C5 w_877_383# a_825_350# 1.88f
C6 w_877_416# p3p2p1g0 1.482f
C7 w_401_n240# b2 1.71f
C8 w_259_n251# p2 1.88f
C9 w_292_n251# a_303_n248# 1.014f
C10 w_802_n14# vdd 1.128f
C11 w_368_n246# b2 1.88f
C12 w_292_n251# a_270_n248# 1.88f
C13 w_259_n251# a_270_n248# 1.014f
C14 w_678_n208# a_615_n203# 1.014f
C15 w_711_68# vdd 1.128f
C16 w_521_464# p2 1.014f
C17 g1 vdd 1.26f
C18 g0 p1p0c0 0.18f
C19 w_602_n213# a_615_n203# 2.82f
C20 w_569_n219# a2 1.014f
C21 w_678_68# vdd 1.128f
C22 w_818_138# c1 1.88f
C23 w_642_625# a_518_635# 1.014f
C24 w_401_n240# a2 1.014f
C25 w_725_411# p2g1 2.312f
C26 w_368_n246# a2 1.17f
C27 w_569_57# vdd 1.128f
C28 w_604_625# a_518_635# 3.59f
C29 g0 p1g0 1.01f
C30 w_504_133# c1 1.88f
C31 w_785_132# a_798_100# 1.88f
C32 w_927_143# a_907_111# 1.014f
C33 a_693_378# gnd 2.424f
C34 w_960_n137# s3 1.88f
C35 w_329_n250# a2 1.128f
C36 w_400_28# vdd 1.128f
C37 w_571_625# a_518_635# 3.59f
C38 w_894_143# a_907_111# 1.88f
C39 w_384_462# p2 1.014f
C40 c3 a_912_n157# 0.54f
C41 w_877_416# a_883_429# 1.41f
C42 w_538_625# a_518_635# 3.59f
C43 w_472_604# a_381_614# 1.014f
C44 w_894_143# a_831_148# 1.014f
C45 w_877_451# a_883_429# 1.41f
C46 w_725_411# a_731_417# 2.444f
C47 w_505_625# a_518_635# 2.45f
C48 w_434_604# a_381_614# 3.59f
C49 w_857_147# a_831_148# 1.128f
C50 w_725_444# a_731_417# 1.128f
C51 w_877_451# p3p2g1 1.482f
C52 w_401_604# a_381_614# 3.59f
C53 w_291_17# vdd 1.128f
C54 w_818_138# a_831_148# 2.162f
C55 w_857_147# a_866_144# 0.936f
C56 w_439_134# a_445_140# 2.444f
C57 w_504_133# a_445_147# 1.014f
C58 b2 a_346_n176# 1.08f
C59 w_725_444# p2p1p0c0 1.482f
C60 w_450_462# g0 1.014f
C61 b0 a_345_92# 1.08f
C62 w_368_604# a_381_614# 2.45f
C63 w_335_599# a_315_567# 1.014f
C64 w_851_n142# c3 1.88f
C65 w_258_17# vdd 1.128f
C66 w_439_134# a_445_147# 1.88f
C67 w_439_167# a_445_140# 1.128f
C68 w_205_450# p2 1.014f
C69 w_857_147# p1 1.128f
C70 w_790_410# a_693_378# 1.014f
C71 w_571_625# p1 1.014f
C72 c1 a_879_123# 0.54f
C73 b0 a_302_20# 6.03f
C74 w_960_n137# a_940_n169# 1.014f
C75 w_302_599# a_315_567# 1.88f
C76 w_226_594# a_206_556# 1.014f
C77 w_927_143# vdd 1.128f
C78 w_642_625# vdd 1.128f
C79 w_818_138# p1 1.17f
C80 b1 gnd 2.314f
C81 b2 a_303_n248# 6.03f
C82 w_725_411# a_693_378# 1.88f
C83 g0 p2 2.07f
C84 w_193_588# a_206_556# 1.88f
C85 w_894_143# vdd 1.128f
C86 a_534_474# p1 0.19f
C87 w_818_n148# a_831_n180# 1.88f
C88 w_927_n137# a_940_n169# 1.88f
C89 w_785_132# p1 1.014f
C90 w_604_625# vdd 1.128f
C91 w_845_654# p3p2p1p0c0 1.88f
C92 w_877_451# a_883_464# 1.598f
C93 b0 a_324_88# 0.54f
C94 a_397_472# p1 0.19f
C95 w_302_599# a_239_604# 1.014f
C96 w_927_n137# a_864_n132# 1.014f
C97 w_571_625# vdd 1.128f
C98 b1 vdd 1.26f
C99 b2 a_325_n180# 0.54f
C100 w_725_444# a_731_457# 1.41f
C101 w_226_594# a_239_604# 2.82f
C102 w_890_n133# a_864_n132# 1.128f
C103 w_258_17# p0 1.88f
C104 a1 vdd 2.52f
C105 w_538_625# vdd 1.128f
C106 w_658_464# p2p1p0c0 1.88f
C107 a0 b0 4.458f
C108 w_851_n142# a_864_n132# 2.162f
C109 w_890_n133# a_899_n136# 0.936f
C110 w_785_132# vdd 1.128f
C111 g0 a_380_291# 1.01f
C112 w_708_654# p2 1.014f
C113 w_505_625# vdd 1.128f
C114 a_612_n65# vdd 1.89f
C115 w_725_479# a_731_457# 1.41f
C116 w_504_133# vdd 1.128f
C117 w_439_167# pocin 1.482f
C118 w_472_604# vdd 1.128f
C119 w_878_485# a_883_464# 1.41f
C120 w_725_479# p2g1g0 1.482f
C121 w_874_1# p2 1.128f
C122 w_400_185# pocin 1.88f
C123 w_434_604# vdd 1.128f
C124 w_878_485# p3g2 1.482f
C125 w_835_n8# p2 1.17f
C126 a_304_328# g0 1.35f
C127 w_439_167# vdd 1.41f
C128 a_534_474# cin 0.19f
C129 w_401_604# vdd 1.128f
C130 a2 b2 3.468f
C131 a_615_73# b0 1.91f
C132 a_534_474# p0 0.19f
C133 w_400_185# vdd 1.128f
C134 w_802_n14# p2 1.014f
C135 w_400_185# a_380_153# 1.014f
C136 w_368_604# vdd 1.128f
C137 a_615_n203# b2 1.91f
C138 w_347_461# p2g1 1.88f
C139 a_251_466# vdd 1.89f
C140 w_708_n70# g1 1.88f
C141 w_367_185# vdd 1.128f
C142 w_367_185# a_380_153# 1.88f
C143 w_291_180# a_271_142# 1.014f
C144 w_505_625# p3 1.014f
C145 w_335_599# vdd 1.128f
C146 w_302_599# vdd 1.128f
C147 w_258_174# a_271_142# 1.88f
C148 w_258_174# vdd 1.128f
C149 w_867_277# vdd 1.128f
C150 w_708_n70# a_688_n102# 1.014f
C151 w_238_456# g1 1.128f
C152 w_193_588# vdd 1.128f
C153 a_864_n132# c3 6.03f
C154 w_834_277# vdd 1.128f
C155 w_675_n70# a_688_n102# 1.88f
C156 w_599_n75# a_579_n113# 1.014f
C157 w_291_180# cin 1.128f
C158 w_368_604# p3 1.014f
C159 w_658_464# a_534_474# 1.014f
C160 w_725_479# a_731_492# 1.598f
C161 w_878_485# a_884_498# 1.598f
C162 w_566_n81# a_579_n113# 1.88f
C163 w_711_68# g0 1.88f
C164 b0 gnd 1.91f
C165 w_620_464# a_534_474# 3.59f
C166 a_831_148# c1 6.03f
C167 w_258_174# p0 1.014f
C168 w_726_513# a_731_492# 1.41f
C169 w_879_518# a_884_498# 1.41f
C170 w_587_464# a_534_474# 3.59f
C171 w_328_n116# a_337_n67# 0.936f
C172 w_725_266# vdd 1.128f
C173 w_367_185# a_304_190# 1.014f
C174 b0 vdd 1.26f
C175 w_554_464# a_534_474# 3.59f
C176 w_488_462# p2p1g0 1.88f
C177 w_400_n106# a_345_n42# 1.88f
C178 w_676_271# vdd 1.128f
C179 w_867_277# s0 1.88f
C180 w_291_180# a_304_190# 2.82f
C181 a0 vdd 2.52f
C182 w_193_588# p3 1.014f
C183 w_521_464# a_534_474# 2.45f
C184 w_758_272# cin 1.88f
C185 w_797_281# p0 1.128f
C186 w_367_n112# a_302_n114# 2.162f
C187 w_758_272# p0 1.17f
C188 w_488_462# a_397_472# 1.014f
C189 a_518_635# p1 0.19f
C190 w_328_n116# a_302_n114# 1.128f
C191 w_611_340# vdd 1.88f
C192 w_725_266# p0 1.014f
C193 w_450_462# a_397_472# 3.59f
C194 w_544_301# vdd 1.128f
C195 w_291_n117# a_302_n114# 1.014f
C196 a_688_664# p1 0.19f
C197 w_440_301# p1 1.014f
C198 a_615_73# vdd 1.89f
C199 a_445_147# gnd 0.808f
C200 w_538_625# p2 1.014f
C201 w_417_462# a_397_472# 3.59f
C202 a_239_604# vdd 1.89f
C203 w_291_n117# a_269_n114# 1.88f
C204 w_599_n75# b1 1.128f
C205 w_506_301# vdd 1.128f
C206 w_725_266# a_738_234# 1.88f
C207 w_384_462# a_397_472# 2.45f
C208 w_473_301# vdd 1.128f
C209 w_258_n117# a_269_n114# 1.014f
C210 w_675_n70# a_612_n65# 1.014f
C211 w_238_456# a_218_418# 1.014f
C212 w_711_n346# g3 1.88f
C213 w_440_301# vdd 1.128f
C214 w_400_n106# b1 1.71f
C215 w_599_n75# a_612_n65# 2.82f
C216 w_566_n81# a1 1.014f
C217 w_226_594# g2 1.128f
C218 w_347_461# a_327_429# 1.014f
C219 w_205_450# a_218_418# 1.88f
C220 w_711_n346# vdd 1.128f
C221 w_604_625# g0 1.014f
C222 w_400_323# vdd 1.128f
C223 w_367_n112# b1 1.88f
C224 w_400_n106# a1 1.014f
C225 w_867_277# a_847_245# 1.014f
C226 w_506_301# cin 1.014f
C227 w_258_312# p1 1.014f
C228 w_401_604# p2 1.014f
C229 w_314_461# a_327_429# 1.88f
C230 w_678_n346# vdd 1.128f
C231 w_367_n112# a1 1.17f
C232 w_367_323# vdd 1.128f
C233 w_944_n3# s2 1.88f
C234 w_834_277# a_847_245# 1.88f
C235 w_328_n116# a1 1.128f
C236 a_688_664# cin 0.19f
C237 w_611_272# p1p0c0 2.312f
C238 w_834_277# a_771_282# 1.014f
C239 w_473_301# p0 1.014f
C240 p1 vdd 2.52f
C241 w_569_n357# vdd 1.128f
C242 w_711_n346# a_691_n378# 1.014f
C243 a_397_472# g0 0.19f
C244 a_688_664# p0 0.19f
C245 w_258_312# vdd 1.128f
C246 w_797_281# a_771_282# 1.128f
C247 w_611_272# a_617_278# 2.444f
C248 w_504_133# g0 1.33f
C249 w_314_461# a_251_466# 1.014f
C250 w_642_625# p3p2p1g0 1.88f
C251 w_678_n346# a_691_n378# 1.88f
C252 w_401_n374# vdd 1.128f
C253 w_602_n351# a_582_n389# 1.014f
C254 w_942_382# vdd 1.128f
C255 w_439_134# g0 2.996f
C256 w_758_272# a_771_282# 2.162f
C257 w_611_305# a_617_278# 1.128f
C258 w_676_271# a_600_239# 1.014f
C259 w_797_281# a_806_278# 0.936f
C260 w_238_456# a_251_466# 2.82f
C261 w_569_n357# a_582_n389# 1.88f
C262 w_835_n8# c2 1.88f
C263 w_544_301# p1p0c0 1.88f
C264 w_611_272# a_600_239# 1.88f
C265 w_611_305# p1g0 1.482f
C266 c2 a_896_n23# 0.54f
C267 w_292_n385# vdd 1.128f
C268 w_329_n384# a_338_n335# 0.936f
C269 w_944_n3# a_924_n35# 1.014f
C270 w_802_n14# a_815_n46# 1.88f
C271 w_259_n385# vdd 1.128f
C272 w_401_n374# a_346_n310# 1.88f
C273 w_790_410# vdd 1.128f
C274 w_911_n3# a_924_n35# 1.88f
C275 cin vdd 1.26f
C276 w_711_n208# vdd 1.128f
C277 w_911_n3# a_848_2# 1.014f
C278 p0 vdd 2.52f
C279 w_678_n208# vdd 1.128f
C280 cin a_819_257# 0.54f
C281 w_874_1# a_848_2# 1.128f
C282 p3 vdd 2.52f
C283 w_611_305# a_617_318# 1.41f
C284 w_602_n351# b3 1.128f
C285 w_368_n380# a_303_n382# 2.162f
C286 w_835_n8# a_848_2# 2.162f
C287 w_874_1# a_883_n2# 0.936f
C288 w_611_340# a_617_318# 1.41f
C289 w_400_323# p1g0 1.88f
C290 w_329_n384# a_303_n382# 1.128f
C291 w_678_n346# a_615_n341# 1.014f
C292 w_569_n219# vdd 1.128f
C293 w_879_518# g3 1.482f
C294 b3 gnd 1.73f
C295 a_304_190# vdd 1.89f
C296 w_401_n240# vdd 1.128f
C297 w_401_n374# b3 1.71f
C298 w_602_n351# a_615_n341# 2.82f
C299 w_259_n385# p3 1.88f
C300 w_569_n357# a3 1.014f
C301 w_292_n385# a_303_n382# 1.014f
C302 w_879_518# vdd 1.88f
C303 w_544_301# a_453_311# 1.014f
C304 w_434_604# g1 1.014f
C305 b1 a_345_n42# 1.08f
C306 w_368_n380# b3 1.88f
C307 w_292_n385# a_270_n382# 1.88f
C308 w_401_n374# a3 1.014f
C309 a_381_614# p2 0.19f
C310 w_726_513# vdd 1.88f
C311 b3 vdd 1.26f
C312 w_506_301# a_453_311# 3.59f
C313 b1 a_302_n114# 6.03f
C314 w_368_n380# a3 1.17f
C315 w_259_n385# a_270_n382# 1.014f
C316 w_658_464# vdd 1.128f
C317 a3 vdd 2.52f
C318 w_473_301# a_453_311# 3.59f
C319 w_554_464# p1 1.014f
C320 a_600_239# gnd 1.616f
C321 w_292_n251# vdd 1.128f
C322 w_329_n384# a3 1.128f
C323 a_518_635# p2 0.19f
C324 w_620_464# vdd 1.128f
C325 a_615_n341# vdd 1.89f
C326 w_440_301# a_453_311# 2.45f
C327 b1 a_324_n46# 0.54f
C328 a_688_664# p2 0.19f
C329 w_259_n251# vdd 1.128f
C330 w_472_604# p3p2g1 1.88f
C331 w_587_464# vdd 1.128f
C332 g0 c1 1.01f
C333 w_960_n137# vdd 1.128f
C334 w_602_63# a_582_25# 1.014f
C335 w_711_68# a_691_36# 1.014f
C336 w_554_464# vdd 1.128f
C337 g2 vdd 1.26f
C338 b3 a_346_n310# 1.08f
C339 w_927_n137# vdd 1.128f
C340 w_675_654# a_688_664# 2.45f
C341 w_678_68# a_691_36# 1.88f
C342 w_569_57# a_582_25# 1.88f
C343 w_521_464# vdd 1.128f
C344 w_417_462# p1 1.014f
C345 w_620_464# cin 1.014f
C346 w_488_462# vdd 1.128f
C347 b3 a_303_n382# 6.03f
C348 a_518_635# g0 0.19f
C349 w_328_18# a_337_67# 0.936f
C350 w_450_462# vdd 1.128f
C351 w_587_464# p0 1.014f
C352 w_400_323# a_380_291# 1.014f
C353 a1 b1 4.008f
C354 w_845_654# a_688_664# 1.014f
C355 g0 a_445_147# 0.72f
C356 w_818_n148# vdd 1.128f
C357 w_711_n208# g2 1.88f
C358 w_417_462# vdd 1.128f
C359 b3 a_325_n314# 0.54f
C360 w_942_382# c4 1.88f
C361 w_367_323# a_380_291# 1.88f
C362 w_291_318# a_271_280# 1.014f
C363 a_612_n65# b1 2.674f
C364 a_848_2# c2 6.03f
C365 w_807_654# a_688_664# 3.59f
C366 a_771_282# cin 6.03f
C367 w_708_n70# vdd 1.128f
C368 w_384_462# vdd 1.128f
C369 w_400_28# a_345_92# 1.88f
C370 p2 vdd 2.52f
C371 w_400_323# g0 1.33f
C372 w_258_312# a_271_280# 1.88f
C373 w_774_654# a_688_664# 3.59f
C374 w_675_n70# vdd 1.128f
C375 w_347_461# vdd 1.128f
C376 a3 b3 3.738f
C377 w_367_323# g0 1.33f
C378 w_877_383# p3p2p1p0c0 2.312f
C379 w_741_654# a_688_664# 3.59f
C380 w_711_n208# a_691_n240# 1.014f
C381 w_890_n133# p3 1.128f
C382 w_602_63# b0 1.128f
C383 w_367_22# a_302_20# 2.162f
C384 w_314_461# vdd 1.128f
C385 w_675_654# vdd 1.128f
C386 a_615_n341# b3 1.91f
C387 b2 gnd 1.91f
C388 w_291_318# g0 1.128f
C389 w_367_323# a_304_328# 1.014f
C390 w_708_654# a_688_664# 3.59f
C391 w_335_599# p3g2 1.88f
C392 a_453_311# cin 0.19f
C393 w_566_n81# vdd 1.128f
C394 w_678_n208# a_691_n240# 1.88f
C395 w_602_n213# a_582_n251# 1.014f
C396 w_851_n142# p3 1.17f
C397 w_328_18# a_302_20# 1.128f
C398 w_291_318# a_304_328# 2.82f
C399 w_818_n148# p3 1.014f
C400 a_453_311# p0 0.19f
C401 w_569_n219# a_582_n251# 1.88f
C402 w_400_n106# vdd 1.128f
C403 w_611_340# g1 1.482f
C404 w_205_450# vdd 1.128f
C405 w_726_513# g2 1.482f
C406 w_400_28# b0 1.71f
C407 w_291_17# a_302_20# 1.014f
C408 w_569_57# a0 1.014f
C409 b2 vdd 1.26f
C410 a_381_614# g1 0.19f
C411 w_258_n117# p1 1.88f
C412 w_845_654# vdd 1.128f
C413 w_367_22# b0 1.88f
C414 w_291_17# a_269_20# 1.88f
C415 w_400_28# a0 1.014f
C416 w_741_654# p1 1.014f
C417 g0 vdd 4.29f
C418 w_329_n250# a_338_n201# 0.936f
C419 w_678_68# a_615_73# 1.014f
C420 w_807_654# vdd 1.128f
C421 w_367_22# a0 1.17f
C422 w_258_17# a_269_20# 1.014f
C423 a_304_328# vdd 1.89f
C424 w_401_n240# a_346_n176# 1.88f
C425 w_291_n117# vdd 1.128f
C426 w_328_18# a0 1.128f
C427 w_602_63# a_615_73# 2.82f
C428 w_774_654# vdd 1.128f
C429 w_675_654# p3 1.014f
C430 w_258_n117# vdd 1.128f
C431 w_741_654# vdd 1.128f
C432 a2 vdd 2.52f
C433 w_944_n3# vdd 1.128f
C434 w_708_654# vdd 1.128f
C435 w_790_410# c3 1.88f
C436 a_615_n203# vdd 1.89f
C437 w_877_383# a_883_389# 2.444f
C438 w_807_654# cin 1.014f
C439 a_825_350# gnd 3.232f
C440 w_602_n213# b2 1.128f
C441 w_368_n246# a_303_n248# 2.162f
C442 w_911_n3# vdd 1.128f
C443 w_676_271# c2 1.88f
C444 gnd 0 1.293863p  
C445 g3 0 65.881004f  
C446 vdd 0 0.952619p  
C447 a_338_n335# 0 3.742f  
C448 a_582_n389# 0 18.082f  
C449 a_691_n378# 0 14.266f  
C450 a_346_n310# 0 14.946f  
C451 p3 0 0.237858p  
C452 a_303_n382# 0 31.139002f  
C453 a_270_n382# 0 14.266f  
C454 a_325_n314# 0 4.916f  
C455 b3 0 85.516f  
C456 a3 0 0.140213p  
C457 a_615_n341# 0 44.863f  
C458 a_912_n157# 0 4.916f  
C459 g2 0 63.907f  
C460 a_338_n201# 0 3.742f  
C461 a_582_n251# 0 18.082f  
C462 a_691_n240# 0 14.266f  
C463 a_346_n176# 0 14.946f  
C464 p2 0 0.28041p  
C465 a_303_n248# 0 31.139002f  
C466 a_270_n248# 0 14.266f  
C467 a_325_n180# 0 4.916f  
C468 b2 0 85.212006f  
C469 s3 0 3.76f  
C470 c3 0 17.83f  
C471 a_831_n180# 0 14.946f  
C472 a2 0 0.137957p  
C473 a_615_n203# 0 44.863f  
C474 a_940_n169# 0 14.266f  
C475 a_864_n132# 0 31.139002f  
C476 a_899_n136# 0 3.742f  
C477 a_896_n23# 0 4.916f  
C478 g1 0 73.370995f  
C479 a_337_n67# 0 3.742f  
C480 a_579_n113# 0 18.082f  
C481 a_688_n102# 0 14.266f  
C482 a_345_n42# 0 14.946f  
C483 a_302_n114# 0 31.139002f  
C484 a_269_n114# 0 14.266f  
C485 a_324_n46# 0 4.916f  
C486 s2 0 3.76f  
C487 c2 0 17.83f  
C488 a_815_n46# 0 14.946f  
C489 b1 0 88.200005f  
C490 a1 0 0.140495p  
C491 a_612_n65# 0 44.863f  
C492 a_924_n35# 0 14.266f  
C493 a_848_2# 0 31.139002f  
C494 a_883_n2# 0 3.742f  
C495 a_337_67# 0 3.742f  
C496 a_582_25# 0 18.082f  
C497 a_879_123# 0 4.916f  
C498 a_691_36# 0 14.266f  
C499 a_345_92# 0 14.946f  
C500 a_302_20# 0 31.139002f  
C501 a_269_20# 0 14.266f  
C502 a_324_88# 0 4.916f  
C503 b0 0 85.82f  
C504 a0 0 0.144276p  
C505 s1 0 3.76f  
C506 c1 0 17.83f  
C507 a_798_100# 0 14.946f  
C508 a_615_73# 0 44.863f  
C509 a_445_140# 0 4.888f  
C510 a_445_147# 0 19.995f  
C511 a_907_111# 0 14.266f  
C512 a_831_148# 0 31.139002f  
C513 a_866_144# 0 3.742f  
C514 p1 0 0.380473p  
C515 pocin 0 28.03f  
C516 a_271_142# 0 18.082f  
C517 a_380_153# 0 14.266f  
C518 a_819_257# 0 4.916f  
C519 a_496_232# 0 1.316f  
C520 cin 0 80.576996f  
C521 p0 0 0.200305p  
C522 s0 0 3.76f  
C523 a_738_234# 0 14.946f  
C524 a_304_190# 0 44.863f  
C525 a_496_251# 0 1.316f  
C526 p1p0c0 0 12.624001f  
C527 a_617_278# 0 4.888f  
C528 p1g0 0 17.794f  
C529 a_600_239# 0 21.439001f  
C530 a_847_245# 0 14.266f  
C531 a_771_282# 0 31.139002f  
C532 a_806_278# 0 3.742f  
C533 a_617_318# 0 2.585f  
C534 a_453_311# 0 17.889f  
C535 c4 0 4.324f  
C536 p3p2p1p0c0 0 12.624001f  
C537 a_271_280# 0 18.082f  
C538 a_380_291# 0 14.266f  
C539 a_610_376# 0 1.316f  
C540 g0 0 0.141479p  
C541 a_304_328# 0 44.863f  
C542 a_440_393# 0 1.316f  
C543 a_610_395# 0 1.316f  
C544 a_883_389# 0 4.888f  
C545 p3p2p1g0 0 18.358f  
C546 a_825_350# 0 23.035f  
C547 p2g1 0 12.06f  
C548 a_610_414# 0 1.316f  
C549 a_440_412# 0 1.316f  
C550 a_731_417# 0 4.888f  
C551 p2p1p0c0 0 18.358f  
C552 a_883_429# 0 2.585f  
C553 p3p2g1 0 30.286f  
C554 a_693_378# 0 22.275f  
C555 a_731_457# 0 2.585f  
C556 p2g1g0 0 25.962f  
C557 a_883_464# 0 2.35f  
C558 p3g2 0 40.25f  
C559 p2p1g0 0 4.324f  
C560 a_218_418# 0 18.082f  
C561 a_534_474# 0 18.744001f  
C562 a_397_472# 0 17.889f  
C563 a_327_429# 0 14.266f  
C564 a_731_492# 0 2.35f  
C565 a_884_498# 0 2.115f  
C566 a_251_466# 0 44.863f  
C567 a_424_535# 0 1.316f  
C568 a_594_537# 0 1.316f  
C569 a_797_547# 0 1.316f  
C570 a_594_556# 0 1.316f  
C571 a_424_554# 0 1.316f  
C572 a_797_566# 0 1.316f  
C573 a_594_575# 0 1.316f  
C574 a_797_585# 0 1.316f  
C575 a_797_604# 0 1.316f  
C576 a_206_556# 0 18.082f  
C577 a_315_567# 0 14.266f  
C578 a_381_614# 0 17.889f  
C579 a_239_604# 0 44.863f  
C580 a_518_635# 0 18.744001f  
C581 a_688_664# 0 19.599f  









 


* * RISING DELAY MEASUREMENT
* Measure the delay for the final carry-out signal (C4)
.measure tran delay_C4 TRIG V(a0) VAL=0.9 RISE=1 TARG V(c4) VAL=0.9 RISE=1

* Measure the delay for each sum signal
.measure tran delay_S0 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s0) VAL=0.9 RISE=1
.measure tran delay_S1 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s1) VAL=0.9 RISE=1
.measure tran delay_S2 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s2) VAL=0.9 RISE=1
.measure tran delay_S3 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s3) VAL=0.9 RISE=1


* FALLING DELAY MEASUREMENT
* Measure the delay for the final carry-out signal (C4)
* .measure tran delay_C4 TRIG V(a0) VAL=0.1 FALL=1 TARG V(c4) VAL=0.1 FALL=1

* * Measure the delay for each sum signal
* .measure tran delay_S0 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s0) VAL=0.1 FALL=1
* .measure tran delay_S1 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s1) VAL=0.1 FALL=1
* .measure tran delay_S2 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s2) VAL=0.1 FALL=1
* .measure tran delay_S3 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s3) VAL=0.1 FALL=1




.control
  set hcopypscolor = 1             
  set color0 = white               
  set color1 = black               
  set color2 = red                 
  set color3 = blue                
  set color4 = coral               
  set color5 = brown    
  set color6 = cyan
  set color7 = chocolate   
  set color8 = chocolate
  set color9 = blueviolet
  set color10 = cadetblue        
  * for testing        
  * tran 1n 160n
  * for delay  
  tran 0.01n 20n 
  * plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+g0 20+g1 22+g2 24+g3   
  * plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+p0 20+p1 22+p2 24+p3                      
  * plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+s0 20+s1 22+s2 24+s3                      
    plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+c4 20+s0 22+s1 24+s2 26+s3  
    plot g3 2+p3g2 4+p3p2g1 6+p3p2p1g0 8+p3p2p1p0c0 10+c4 
  * plot s0 2+s1 4+s2 6+s3    
        
.endc
