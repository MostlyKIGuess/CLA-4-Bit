* SPICE3 file created from cla.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={40*LAMBDA}
.param width_N={20*LAMBDA}
.global gnd vdd

* Power Supply for the circuit
Vdd vdd gnd 'SUPPLY'


* Input Signals
* for testing
* Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
* Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 30n 60n)     
* Va1 a1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 10n 20n)    
* Vb1 b1 gnd PULSE(0 'SUPPLY' 5n 0.01n 0.01n 30n 60n)    
* Va2 a2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 10n 20n)   
* Vb2 b2 gnd PULSE(0 'SUPPLY' 10n 0.01n 0.01n 30n 60n)   
* Va3 a3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 10n 20n)   
* Vb3 b3 gnd PULSE(0 'SUPPLY' 15n 0.01n 0.01n 30n 60n)   
* Vcin cin gnd DC 0         

* Input Signals for delay measurement
*  rising
Vclk clk gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)  
Va0 a0 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)     
Vb0 b0 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)     
Va1 a1 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)    
Vb1 b1 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)    
Va2 a2 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Vb2 b2 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Va3 a3 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Vb3 b3 gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)   
Vcin cin gnd PULSE(0 'SUPPLY' 10ns 0.01n 0.01n 10n 20n)


* Input Signals for delay measurement
*  falling
* Vclk clk gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)  
* Va0 a0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Vb0 b0 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)     
* Va1 a1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
* Vb1 b1 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)    
* Va2 a2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Vb2 b2 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Va3 a3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Vb3 b3 gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)   
* Vcin cin gnd PULSE(0 'SUPPLY' 0 0.01n 0.01n 10n 20n)                             





* SPICE3 file created from testing.ext - technology: scmos

.option scale=0.09u

M1000 a_445_147# g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 a_691_n240# a_615_n203# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1002 a_615_n203# a_582_n251# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 p2g1 a_327_429# vdd w_347_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_594_575# p1 a_594_556# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1005 a_440_412# p1 a_440_393# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1006 p1p0c0 a_453_311# vdd w_544_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1007 a3 b3 a_303_n382# w_329_n384# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1008 a_848_2# p2 c2 w_835_n8# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1009 a_518_635# p3 vdd w_505_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1010 a_731_457# p2p1p0c0 a_731_417# w_725_444# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1011 b2 a2 a_303_n248# w_368_n246# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1012 gnd a_303_n248# a_270_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1013 p3p2g1 a_381_614# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 p2p1p0c0 a_534_474# vdd w_658_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1015 a_610_395# p1 a_610_377# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1016 b2 a_325_n180# a_303_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1017 a_815_n46# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1018 a_518_635# g0 a_594_575# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1019 a_940_n169# a_864_n132# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1020 s2 a_924_n35# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1021 vdd a0 a_324_88# w_400_28# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 vdd a_302_20# a_269_20# w_291_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1023 a_325_n180# b2 a_303_n248# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1024 g0 a_691_36# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1025 a_825_350# p3p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1026 a_847_245# a_771_282# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 a_304_190# a_271_142# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1028 a_884_498# p3g2 a_883_464# w_878_485# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1029 g3 a_691_n378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 a_731_492# p2p1g0 a_731_457# w_725_479# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1031 a_831_148# a_798_100# c1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1032 a_615_n341# a3 b3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1033 a_831_148# c1 p1 w_857_146# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1034 a_798_100# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1035 a_315_567# a_239_604# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1036 g2 a_691_n240# vdd w_711_n208# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1037 a_582_n251# a2 vdd w_569_n219# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1038 p3g2 a_315_567# vdd w_335_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1039 vdd g3 a_884_498# w_879_518# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1040 a_825_350# p3p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1041 pocin a_380_153# vdd w_400_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1042 vdd a_269_20# p0 w_258_17# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1043 a_218_418# p2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1044 a_380_153# a_304_190# vdd w_367_185# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1045 b1 a1 a_302_n114# w_367_n112# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1046 a_691_36# a_615_73# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1047 a_825_350# p3p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1048 a_271_280# p1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1049 a_907_111# a_831_148# vdd w_894_143# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1050 s2 a_924_n35# vdd w_944_n3# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1051 p3p2p1g0 a_518_635# vdd w_642_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1052 a_615_n203# a_582_n251# b2 w_602_n213# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1053 a_239_604# a_206_556# g2 w_226_594# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1054 a_304_190# a_271_142# cin w_291_180# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1055 a_612_n65# a_579_n113# b1 w_599_n75# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_582_25# a0 vdd w_569_57# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1057 p2p1g0 a_397_472# vdd w_488_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 c3 a_693_378# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1059 a_440_393# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1060 a_612_n65# a_579_n113# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1061 a_924_n35# a_848_2# vdd w_911_n3# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1062 a_688_664# p0 vdd w_774_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 a_445_147# pocin gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1064 p2g1 a_327_429# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1065 a_600_239# p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1066 s3 a_940_n169# vdd w_960_n137# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1067 a_327_429# a_251_466# vdd w_314_461# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1068 a_848_2# a_815_n46# c2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1069 a_688_664# cin vdd w_807_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1070 a_693_378# p2g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1071 a_251_466# p2 g1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1072 a_325_n314# b3 a_303_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1073 a_688_n102# a_612_n65# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1074 a_738_234# p0 vdd w_725_266# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_924_n35# a_848_2# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1076 p3p2g1 a_381_614# vdd w_472_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1077 a_206_556# p3 vdd w_193_588# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1078 a_424_535# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1079 g2 a_691_n240# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1080 a_610_377# p2 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1081 s0 a_847_245# vdd w_867_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1082 a_582_n389# a3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1083 a_691_n378# a_615_n341# vdd w_678_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1084 a_864_n132# a_831_n180# c3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1085 vdd a2 a_325_n180# w_401_n240# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1086 a_615_n203# a2 b2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1087 g1 a_688_n102# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1088 c4 a_825_350# vdd w_942_382# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1089 a_424_554# p2 a_424_535# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1090 a_453_311# p0 vdd w_473_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1091 a_831_n180# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1092 a_315_567# a_239_604# vdd w_302_599# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1093 p3p2p1p0c0 a_688_664# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1094 a_771_282# p0 cin w_758_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1095 a_271_142# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1096 a_612_n65# a1 b1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1097 a_534_474# cin vdd w_620_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1098 a_534_474# p0 vdd w_587_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1099 a_453_311# cin vdd w_506_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1100 a_271_280# p1 vdd w_258_312# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1101 a_693_378# p2p1g0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1102 a_381_614# g1 a_424_554# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1103 a_883_429# p3p2p1g0 a_883_389# w_877_416# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1104 c1 a_445_147# vdd w_504_133# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1105 a_304_328# a_271_280# g0 w_291_318# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1106 a_825_350# p3g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1107 a_688_664# p1 vdd w_741_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1108 a_797_604# p0 a_797_585# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1109 vdd a_269_n114# p1 w_258_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1110 p1g0 a_380_291# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1111 a_324_n46# b1 a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_327_429# a_251_466# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1113 a1 b1 a_302_n114# w_328_n116# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1114 s1 a_907_111# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1115 a_693_378# p2p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1116 a_380_291# a_304_328# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1117 c2 a_600_239# vdd w_676_271# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1118 b0 a_324_88# a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1119 b3 a3 a_303_n382# w_368_n380# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1120 a_688_n102# a_612_n65# vdd w_675_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 b1 a_324_n46# a_302_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1122 a_815_n46# p2 vdd w_802_n14# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 vdd a3 a_325_n314# w_401_n374# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1124 a_615_73# a_582_25# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1125 p1p0c0 a_453_311# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1126 a_324_88# b0 a_302_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1127 a_688_664# cin a_797_604# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1128 vdd g2 a_731_492# w_726_513# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1129 a_883_464# p3p2g1 a_883_429# w_877_451# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1130 a_693_378# g2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1131 g1 a_688_n102# vdd w_708_n70# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1132 a_831_148# c1 a_798_100# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 a_864_n132# p3 c3 w_851_n142# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1134 a_304_328# p1 g0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1135 a_771_282# a_738_234# cin Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1136 a_518_635# p1 vdd w_571_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1137 a_397_472# g0 vdd w_450_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1138 a_579_n113# a1 vdd w_566_n81# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1139 a_797_547# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1140 a_496_251# p0 a_496_232# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1141 a_848_2# c2 p2 w_874_0# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1142 a_518_635# g0 vdd w_604_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1143 a_825_350# p3p2p1p0c0 a_883_389# w_877_383# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1144 p2p1p0c0 a_534_474# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1145 g0 a_691_36# vdd w_711_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1146 a_847_245# a_771_282# vdd w_834_277# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1147 vdd a_270_n248# p2 w_259_n251# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1148 a_579_n113# a1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1149 a_239_604# a_206_556# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1150 a_797_566# p2 a_797_547# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1151 a_453_311# cin a_496_251# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1152 a_453_311# p1 vdd w_440_301# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1153 a_798_100# p1 vdd w_785_132# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1154 gnd a3 a_325_n314# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1155 a_534_474# p1 vdd w_554_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1156 a_304_328# a_271_280# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1157 a_445_147# g0 a_445_140# w_439_134# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1158 a_940_n169# a_864_n132# vdd w_927_n137# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1159 a_797_585# p1 a_797_566# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1160 a_864_n132# c3 a_831_n180# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1161 gnd a_302_n114# a_269_n114# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1162 a_691_36# a_615_73# vdd w_678_68# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1163 s3 a_940_n169# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1164 a_864_n132# c3 p3 w_890_n134# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1165 gnd a_269_n114# p1 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1166 a_381_614# g1 vdd w_434_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1167 vdd a_303_n248# a_270_n248# w_292_n251# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1168 pocin a_380_153# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1169 a_848_2# c2 a_815_n46# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1170 a_380_153# a_304_190# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1171 a_831_148# p1 c1 w_818_138# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1172 a_688_664# p3 vdd w_675_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1173 g3 a_691_n378# vdd w_711_n346# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1174 a_907_111# a_831_148# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1175 p1g0 a_380_291# vdd w_400_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1176 c2 a_600_239# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1177 a_615_73# a0 b0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1178 a0 b0 a_302_20# w_328_18# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1179 a_380_291# a_304_328# vdd w_367_323# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1180 vdd a_270_n382# p3 w_259_n385# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1181 a_582_25# a0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1182 a_688_664# p2 vdd w_708_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1183 p2p1g0 a_397_472# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1184 gnd a2 a_325_n180# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1185 vdd pocin a_445_140# w_439_167# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 c3 a_693_378# vdd w_790_410# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1187 a_304_190# p0 cin Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1188 a_251_466# a_218_418# g1 w_238_456# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1189 vdd a1 a_324_n46# w_400_n106# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1190 a_397_472# g0 a_440_412# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1191 a_691_n378# a_615_n341# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1192 a_615_n341# a_582_n389# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1193 a_397_472# p2 vdd w_384_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1194 vdd a_303_n382# a_270_n382# w_292_n385# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1195 vdd a_302_n114# a_269_n114# w_291_n117# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1196 a_617_318# p1g0 a_617_278# w_611_305# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1197 a_771_282# cin p0 w_797_280# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1198 a_738_234# p0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1199 a_691_n240# a_615_n203# vdd w_678_n208# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1200 a_518_635# p2 vdd w_538_625# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1201 a_496_232# p1 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1202 b0 a0 a_302_20# w_367_22# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1203 a_397_472# p1 vdd w_417_462# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_206_556# p3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1205 gnd a_270_n382# p3 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1206 a_610_414# p0 a_610_395# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1207 p3p2p1p0c0 a_688_664# vdd w_845_654# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1208 a_271_142# p0 vdd w_258_174# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1209 a_582_n251# a2 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1210 a_534_474# p2 vdd w_521_464# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1211 s0 a_847_245# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1212 vdd g1 a_617_318# w_611_340# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1213 c4 a_825_350# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 gnd a0 a_324_88# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1215 gnd a1 a_324_n46# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1216 gnd a_302_20# a_269_20# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1217 a_381_614# p2 vdd w_401_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1218 a_534_474# cin a_610_414# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1219 a2 b2 a_303_n248# w_329_n250# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1220 a_251_466# a_218_418# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1221 a_771_282# cin a_738_234# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1222 a_381_614# p3 vdd w_368_604# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1223 p3g2 a_315_567# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1224 a_594_537# p3 gnd Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1225 a_600_239# g1 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1226 a_615_73# a_582_25# b0 w_602_63# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1227 a_582_n389# a3 vdd w_569_n357# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1228 a_239_604# p3 g2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1229 b3 a_325_n314# a_303_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1230 gnd a_303_n382# a_270_n382# Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1231 a_218_418# p2 vdd w_205_450# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1232 a_825_350# g3 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1233 a_600_239# p1p0c0 a_617_278# w_611_272# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1234 s1 a_907_111# vdd w_927_143# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1235 c1 a_445_147# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1236 p3p2p1g0 a_518_635# gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1237 a_693_378# p2g1 a_731_417# w_725_411# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1238 a_831_n180# p3 vdd w_818_n148# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1239 a_600_239# p1p0c0 gnd Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1240 gnd a_270_n248# p2 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1241 a_594_556# p2 a_594_537# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1242 gnd a_269_20# p0 Gnd CMOSN w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1243 a_615_n341# a_582_n389# b3 w_602_n351# CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
C0 w_400_323# g0 1.33f
C1 w_942_382# c4 1.88f
C2 b1 a_302_n114# 4.68f
C3 w_774_654# a_688_664# 3.59f
C4 w_292_n385# vdd 1.128f
C5 g0 a_445_147# 0.72f
C6 w_367_323# g0 1.33f
C7 w_741_654# a_688_664# 3.59f
C8 w_259_n385# vdd 1.128f
C9 w_602_n351# b3 1.128f
C10 w_368_n380# a_303_n382# 2.162f
C11 w_790_410# vdd 1.128f
C12 w_291_318# g0 1.128f
C13 w_877_383# p3p2p1p0c0 2.202f
C14 w_367_323# a_304_328# 1.014f
C15 cin vdd 1.26f
C16 b1 a_324_n46# 2.925f
C17 w_708_654# a_688_664# 3.59f
C18 w_401_n374# a_325_n314# 1.88f
C19 w_329_n384# a_303_n382# 1.128f
C20 w_678_n346# a_615_n341# 1.014f
C21 a_453_311# cin 0.19f
C22 w_711_n208# vdd 1.128f
C23 w_291_318# a_304_328# 2.82f
C24 p0 vdd 2.52f
C25 w_401_n374# b3 1.71f
C26 w_602_n351# a_615_n341# 2.82f
C27 w_569_n357# a3 1.014f
C28 w_292_n385# a_303_n382# 1.014f
C29 a_453_311# p0 0.19f
C30 w_678_n208# vdd 1.128f
C31 w_602_63# b0 1.128f
C32 w_367_22# a_302_20# 2.162f
C33 w_368_n380# b3 1.88f
C34 w_292_n385# a_270_n382# 1.88f
C35 w_401_n374# a3 1.014f
C36 w_400_28# a_324_88# 1.88f
C37 w_328_18# a_302_20# 1.128f
C38 w_642_625# vdd 1.128f
C39 w_569_n219# vdd 1.128f
C40 w_368_n380# a3 1.17f
C41 w_329_n384# b3 1.17f
C42 w_259_n385# a_270_n382# 1.014f
C43 w_258_n117# p1 1.88f
C44 w_400_28# b0 1.71f
C45 w_291_17# a_302_20# 1.014f
C46 w_569_57# a0 1.014f
C47 w_879_518# g3 1.482f
C48 w_741_654# p1 1.014f
C49 a_304_190# vdd 1.89f
C50 a1 b1 4.008f
C51 w_604_625# vdd 1.128f
C52 w_329_n384# a3 1.128f
C53 w_401_n240# vdd 1.128f
C54 w_367_22# b0 1.88f
C55 w_291_17# a_269_20# 1.88f
C56 w_400_28# a0 1.014f
C57 w_678_68# a_615_73# 1.014f
C58 w_879_518# vdd 1.88f
C59 a_612_n65# b1 2.674f
C60 w_571_625# vdd 1.128f
C61 w_367_22# a0 1.17f
C62 w_328_18# b0 1.17f
C63 w_258_17# a_269_20# 1.014f
C64 w_726_513# vdd 1.88f
C65 w_602_63# a_615_73# 2.82f
C66 w_538_625# vdd 1.128f
C67 w_328_18# a0 1.128f
C68 w_658_464# vdd 1.128f
C69 w_807_654# cin 1.014f
C70 w_877_383# a_883_389# 2.444f
C71 a_600_239# gnd 1.616f
C72 c2 a_815_n46# 1.845f
C73 w_505_625# vdd 1.128f
C74 w_292_n251# vdd 1.128f
C75 w_620_464# vdd 1.128f
C76 w_877_416# a_883_389# 1.128f
C77 w_942_382# a_825_350# 1.014f
C78 w_472_604# vdd 1.128f
C79 w_259_n251# vdd 1.128f
C80 w_434_604# g1 1.014f
C81 w_587_464# vdd 1.128f
C82 w_774_654# p0 1.014f
C83 w_877_383# a_825_350# 1.88f
C84 w_877_416# p3p2p1g0 1.482f
C85 w_434_604# vdd 1.128f
C86 w_960_n137# vdd 1.128f
C87 w_554_464# vdd 1.128f
C88 w_401_604# vdd 1.128f
C89 w_927_n137# vdd 1.128f
C90 w_711_n208# a_691_n240# 1.014f
C91 w_604_625# g0 1.014f
C92 w_521_464# vdd 1.128f
C93 w_927_143# s1 1.88f
C94 g1 gnd 15.03f
C95 w_368_604# vdd 1.128f
C96 w_678_n208# a_691_n240# 1.88f
C97 w_602_n213# a_582_n251# 1.014f
C98 w_488_462# vdd 1.128f
C99 c2 a_848_2# 4.68f
C100 w_335_599# vdd 1.128f
C101 g0 p1p0c0 0.18f
C102 w_569_n219# a_582_n251# 1.88f
C103 w_450_462# vdd 1.128f
C104 g1 vdd 2.472f
C105 w_302_599# vdd 1.128f
C106 w_818_n148# vdd 1.128f
C107 w_417_462# vdd 1.128f
C108 w_708_n70# g1 1.88f
C109 w_725_411# p2g1 2.202f
C110 w_708_n70# vdd 1.128f
C111 g0 p1g0 1.01f
C112 w_642_625# p3p2p1g0 1.88f
C113 w_384_462# vdd 1.128f
C114 w_193_588# vdd 1.128f
C115 w_675_n70# vdd 1.128f
C116 a_206_556# g2 0.846f
C117 w_857_146# c1 1.17f
C118 w_347_461# vdd 1.128f
C119 w_785_132# a_798_100# 1.88f
C120 w_877_416# a_883_429# 1.41f
C121 w_602_n213# b2 1.128f
C122 w_368_n246# a_303_n248# 2.162f
C123 w_927_143# a_907_111# 1.014f
C124 w_818_138# c1 1.88f
C125 w_314_461# vdd 1.128f
C126 w_675_654# vdd 1.128f
C127 w_238_456# g1 2.724f
C128 w_877_451# a_883_429# 1.41f
C129 w_725_411# a_731_417# 2.444f
C130 w_401_n240# a_325_n180# 1.88f
C131 w_329_n250# a_303_n248# 1.128f
C132 w_566_n81# vdd 1.128f
C133 w_894_143# a_907_111# 1.88f
C134 b3 gnd 1.73f
C135 w_205_450# g1 1.596f
C136 w_725_444# a_731_417# 1.128f
C137 w_877_451# p3p2g1 1.482f
C138 w_400_n106# vdd 1.128f
C139 w_401_n240# b2 1.71f
C140 w_292_n251# a_303_n248# 1.014f
C141 w_894_143# a_831_148# 1.014f
C142 w_205_450# vdd 1.128f
C143 w_504_133# c1 1.88f
C144 w_676_271# c2 1.88f
C145 a_239_604# g2 0.786f
C146 w_725_444# p2p1p0c0 1.482f
C147 w_450_462# g0 1.014f
C148 w_368_n246# b2 1.88f
C149 w_292_n251# a_270_n248# 1.88f
C150 w_678_n208# a_615_n203# 1.014f
C151 w_857_146# a_831_148# 1.128f
C152 w_845_654# vdd 1.128f
C153 b3 vdd 0.72f
C154 w_790_410# a_693_378# 1.014f
C155 g0 vdd 4.29f
C156 w_602_n213# a_615_n203# 2.82f
C157 w_569_n219# a2 1.014f
C158 w_329_n250# b2 1.17f
C159 w_259_n251# a_270_n248# 1.014f
C160 w_439_134# a_445_140# 2.444f
C161 w_504_133# a_445_147# 1.014f
C162 w_818_138# a_831_148# 2.162f
C163 w_807_654# vdd 1.128f
C164 w_857_146# p1 1.128f
C165 w_790_410# c3 1.88f
C166 a3 vdd 2.52f
C167 w_725_411# a_693_378# 1.88f
C168 a_304_328# vdd 1.89f
C169 w_291_n117# vdd 1.128f
C170 a_534_474# p1 0.19f
C171 w_401_n240# a2 1.014f
C172 w_259_n385# p3 1.88f
C173 w_818_138# p1 1.17f
C174 w_439_134# a_445_147# 1.88f
C175 w_439_167# a_445_140# 1.128f
C176 w_774_654# vdd 1.128f
C177 a_615_n341# vdd 1.08f
C178 w_877_451# a_883_464# 1.598f
C179 a_397_472# p1 0.19f
C180 w_258_n117# vdd 1.128f
C181 w_368_n246# a2 1.17f
C182 w_741_654# vdd 1.128f
C183 w_785_132# p1 1.014f
C184 b3 a_303_n382# 4.68f
C185 w_725_444# a_731_457# 1.41f
C186 w_845_654# p3p2p1p0c0 1.88f
C187 a_381_614# p2 0.19f
C188 w_944_n3# vdd 1.128f
C189 w_329_n250# a2 1.128f
C190 w_258_17# p0 1.88f
C191 w_708_654# vdd 1.128f
C192 w_658_464# p2p1p0c0 1.88f
C193 a_825_350# gnd 3.232f
C194 b0 a_302_20# 4.68f
C195 g0 a_380_291# 1.01f
C196 w_960_n137# s3 1.88f
C197 w_911_n3# vdd 1.128f
C198 b3 a_325_n314# 2.925f
C199 w_725_479# a_731_457# 1.41f
C200 a_518_635# p2 0.19f
C201 b2 gnd 1.91f
C202 w_878_485# a_883_464# 1.41f
C203 w_725_479# p2p1g0 1.482f
C204 b0 a_324_88# 2.925f
C205 a_688_664# p2 0.19f
C206 a_534_474# cin 0.19f
C207 w_439_167# pocin 1.482f
C208 a3 b3 3.738f
C209 w_878_485# p3g2 1.482f
C210 a_304_328# g0 1.35f
C211 w_802_n14# vdd 1.128f
C212 a_534_474# p0 0.19f
C213 w_472_604# p3p2g1 1.88f
C214 w_400_185# pocin 1.88f
C215 b2 vdd 0.9f
C216 a_615_n341# b3 1.91f
C217 a0 b0 4.458f
C218 w_711_68# vdd 1.128f
C219 w_960_n137# a_940_n169# 1.014f
C220 w_347_461# p2g1 1.88f
C221 w_505_625# p3 1.014f
C222 w_678_68# vdd 1.128f
C223 w_818_n148# a_831_n180# 1.88f
C224 w_927_n137# a_940_n169# 1.88f
C225 w_400_185# a_380_153# 1.014f
C226 w_927_n137# a_864_n132# 1.014f
C227 w_367_185# a_380_153# 1.88f
C228 w_291_180# a_271_142# 1.014f
C229 w_711_n208# g2 1.88f
C230 a2 vdd 2.52f
C231 g1 a_615_n203# 2.97f
C232 a_615_73# b0 1.91f
C233 w_890_n134# a_864_n132# 1.128f
C234 w_569_57# vdd 1.128f
C235 w_258_174# a_271_142# 1.88f
C236 a_615_n203# vdd 1.35f
C237 a_693_378# gnd 2.424f
C238 w_400_28# vdd 1.128f
C239 w_851_n142# a_864_n132# 2.162f
C240 w_890_n134# c3 1.17f
C241 w_725_479# a_731_492# 1.598f
C242 w_658_464# a_534_474# 1.014f
C243 w_368_604# p3 1.014f
C244 w_851_n142# c3 1.88f
C245 w_890_n134# p3 1.128f
C246 w_291_180# cin 1.128f
C247 w_878_485# a_884_498# 1.598f
C248 w_488_462# p2p1g0 1.88f
C249 w_620_464# a_534_474# 3.59f
C250 w_851_n142# p3 1.17f
C251 w_711_68# g0 1.88f
C252 w_726_513# a_731_492# 1.41f
C253 w_587_464# a_534_474# 3.59f
C254 c1 a_798_100# 1.845f
C255 g1 p3 83.43f
C256 w_291_17# vdd 1.128f
C257 w_818_n148# p3 1.014f
C258 w_258_174# p0 1.014f
C259 p3 vdd 2.52f
C260 w_554_464# a_534_474# 3.59f
C261 w_879_518# a_884_498# 1.41f
C262 w_726_513# g2 1.482f
C263 w_258_17# vdd 1.128f
C264 w_335_599# p3g2 1.88f
C265 w_367_185# a_304_190# 1.014f
C266 w_521_464# a_534_474# 2.45f
C267 w_193_588# p3 1.014f
C268 w_927_143# vdd 1.128f
C269 w_797_280# cin 1.17f
C270 w_867_277# s0 1.88f
C271 w_291_180# a_304_190# 2.82f
C272 w_894_143# vdd 1.128f
C273 a_218_418# g1 1.212f
C274 w_708_n70# a_688_n102# 1.014f
C275 w_758_272# cin 1.88f
C276 w_797_280# p0 1.128f
C277 b2 a_303_n248# 4.68f
C278 w_675_654# p3 1.014f
C279 w_488_462# a_397_472# 1.014f
C280 w_675_n70# a_688_n102# 1.88f
C281 w_599_n75# a_579_n113# 1.014f
C282 w_758_272# p0 1.17f
C283 w_450_462# a_397_472# 3.59f
C284 w_566_n81# a_579_n113# 1.88f
C285 w_725_266# p0 1.014f
C286 b2 a_325_n180# 2.925f
C287 w_417_462# a_397_472# 3.59f
C288 a_831_148# c1 4.68f
C289 a_518_635# p1 0.19f
C290 w_785_132# vdd 1.128f
C291 b1 gnd 2.314f
C292 w_384_462# a_397_472# 2.45f
C293 g2 gnd 30.06f
C294 w_538_625# p2 1.014f
C295 w_504_133# vdd 1.128f
C296 a_688_664# p1 0.19f
C297 w_725_266# a_738_234# 1.88f
C298 w_440_301# p1 1.014f
C299 w_238_456# a_218_418# 1.014f
C300 b1 vdd 0.9f
C301 w_347_461# a_327_429# 1.014f
C302 w_205_450# a_218_418# 1.88f
C303 g1 a1 16.199999f
C304 g2 vdd 2.068f
C305 w_439_167# vdd 1.41f
C306 w_367_n112# a_302_n114# 2.162f
C307 w_259_n251# p2 1.88f
C308 w_226_594# g2 2.268f
C309 a1 vdd 2.52f
C310 a2 b2 3.468f
C311 w_314_461# a_327_429# 1.88f
C312 a_251_466# g1 1.212f
C313 w_400_n106# a_324_n46# 1.88f
C314 w_328_n116# a_302_n114# 1.128f
C315 w_400_185# vdd 1.128f
C316 w_193_588# g2 1.064f
C317 w_867_277# a_847_245# 1.014f
C318 w_506_301# cin 1.014f
C319 a_615_n203# b2 1.91f
C320 a_612_n65# vdd 1.35f
C321 a_251_466# vdd 1.89f
C322 w_401_604# p2 1.014f
C323 w_291_n117# a_302_n114# 1.014f
C324 w_367_185# vdd 1.128f
C325 w_599_n75# b1 1.128f
C326 w_258_312# p1 1.014f
C327 w_834_277# a_847_245# 1.88f
C328 w_521_464# p2 1.014f
C329 a_397_472# g0 0.19f
C330 w_291_n117# a_269_n114# 1.88f
C331 a_688_664# cin 0.19f
C332 w_675_n70# a_612_n65# 1.014f
C333 w_611_272# p1p0c0 2.202f
C334 w_473_301# p0 1.014f
C335 w_834_277# a_771_282# 1.014f
C336 w_258_n117# a_269_n114# 1.014f
C337 w_258_174# vdd 1.128f
C338 a_688_664# p0 0.19f
C339 w_400_n106# b1 1.71f
C340 w_599_n75# a_612_n65# 2.82f
C341 w_566_n81# a1 1.014f
C342 w_504_133# g0 1.33f
C343 w_797_280# a_771_282# 1.128f
C344 w_611_272# a_617_278# 2.444f
C345 w_314_461# a_251_466# 1.014f
C346 g1 p2 3.825f
C347 w_867_277# vdd 1.128f
C348 w_367_n112# b1 1.88f
C349 w_400_n106# a1 1.014f
C350 w_642_625# a_518_635# 1.014f
C351 w_758_272# a_771_282# 2.162f
C352 w_611_305# a_617_278# 1.128f
C353 w_676_271# a_600_239# 1.014f
C354 w_439_134# g0 2.943f
C355 p2 vdd 2.52f
C356 w_238_456# a_251_466# 2.82f
C357 w_834_277# vdd 1.128f
C358 w_367_n112# a1 1.17f
C359 w_328_n116# b1 1.17f
C360 w_604_625# a_518_635# 3.59f
C361 w_611_272# a_600_239# 1.88f
C362 w_611_305# p1g0 1.482f
C363 w_384_462# p2 1.014f
C364 w_544_301# p1p0c0 1.88f
C365 c3 a_831_n180# 1.845f
C366 w_944_n3# s2 1.88f
C367 w_328_n116# a1 1.128f
C368 w_571_625# a_518_635# 3.59f
C369 g2 a_615_n341# 1.485f
C370 w_472_604# a_381_614# 1.014f
C371 w_538_625# a_518_635# 3.59f
C372 w_725_266# vdd 1.128f
C373 w_505_625# a_518_635# 2.45f
C374 w_434_604# a_381_614# 3.59f
C375 b0 gnd 1.91f
C376 w_676_271# vdd 1.128f
C377 w_401_604# a_381_614# 3.59f
C378 w_611_305# a_617_318# 1.41f
C379 w_205_450# p2 1.014f
C380 c3 a_864_n132# 4.68f
C381 w_368_604# a_381_614# 2.45f
C382 w_335_599# a_315_567# 1.014f
C383 w_611_340# a_617_318# 1.41f
C384 b0 vdd 0.9f
C385 w_802_n14# a_815_n46# 1.88f
C386 w_944_n3# a_924_n35# 1.014f
C387 w_302_599# a_315_567# 1.88f
C388 w_226_594# a_206_556# 1.014f
C389 w_611_340# g1 1.482f
C390 w_400_323# p1g0 1.88f
C391 a0 vdd 2.52f
C392 w_571_625# p1 1.014f
C393 w_611_340# vdd 1.88f
C394 a_381_614# g1 0.19f
C395 w_911_n3# a_924_n35# 1.88f
C396 w_193_588# a_206_556# 1.88f
C397 w_911_n3# a_848_2# 1.014f
C398 w_544_301# vdd 1.128f
C399 w_302_599# a_239_604# 1.014f
C400 w_544_301# a_453_311# 1.014f
C401 a_239_604# vdd 1.89f
C402 w_874_0# a_848_2# 1.128f
C403 w_506_301# vdd 1.128f
C404 w_226_594# a_239_604# 2.82f
C405 w_506_301# a_453_311# 3.59f
C406 w_708_654# p2 1.014f
C407 a_615_73# vdd 1.35f
C408 a_738_234# cin 1.845f
C409 w_835_n8# a_848_2# 2.162f
C410 w_874_0# c2 1.17f
C411 w_473_301# vdd 1.128f
C412 w_473_301# a_453_311# 3.59f
C413 a_445_147# gnd 0.808f
C414 w_711_n346# g3 1.88f
C415 w_835_n8# c2 1.88f
C416 w_874_0# p2 1.128f
C417 w_440_301# vdd 1.128f
C418 w_440_301# a_453_311# 2.45f
C419 w_554_464# p1 1.014f
C420 w_711_n346# vdd 1.128f
C421 w_400_323# vdd 1.128f
C422 w_835_n8# p2 1.17f
C423 w_678_n346# vdd 1.128f
C424 w_802_n14# p2 1.014f
C425 w_367_323# vdd 1.128f
C426 w_675_654# a_688_664# 2.45f
C427 w_711_n346# a_691_n378# 1.014f
C428 w_620_464# cin 1.014f
C429 w_569_n357# vdd 1.128f
C430 w_678_n346# a_691_n378# 1.88f
C431 w_602_n351# a_582_n389# 1.014f
C432 w_258_312# vdd 1.128f
C433 w_417_462# p1 1.014f
C434 w_291_318# a_271_280# 1.014f
C435 p1 vdd 2.52f
C436 g2 p3 1.575f
C437 w_569_n357# a_582_n389# 1.88f
C438 w_401_n374# vdd 1.128f
C439 a_518_635# g0 0.19f
C440 w_942_382# vdd 1.128f
C441 w_711_68# a_691_36# 1.014f
C442 w_587_464# p0 1.014f
C443 w_258_312# a_271_280# 1.88f
C444 w_400_323# a_380_291# 1.014f
C445 w_845_654# a_688_664# 1.014f
C446 g0 c1 1.01f
C447 w_678_68# a_691_36# 1.88f
C448 w_602_63# a_582_25# 1.014f
C449 w_367_323# a_380_291# 1.88f
C450 w_807_654# a_688_664# 3.59f
C451 a_771_282# cin 4.68f
C452 w_569_57# a_582_25# 1.88f
C453 gnd 0 1.283899p  
C454 g3 0 65.881004f  
C455 vdd 0 0.955556p  
C456 a_582_n389# 0 18.082f  
C457 a_691_n378# 0 14.266f  
C458 a_303_n382# 0 30.763f  
C459 a_270_n382# 0 14.266f  
C460 a_325_n314# 0 26.066f  
C461 b3 0 90.43f  
C462 a3 0 0.140213p  
C463 a_615_n341# 0 44.863f  
C464 a_582_n251# 0 18.082f  
C465 a_691_n240# 0 14.266f  
C466 a_303_n248# 0 30.763f  
C467 a_270_n248# 0 14.266f  
C468 a_325_n180# 0 26.066f  
C469 b2 0 90.126f  
C470 s3 0 3.76f  
C471 a_831_n180# 0 26.066f  
C472 a2 0 0.137957p  
C473 a_615_n203# 0 44.863f  
C474 a_940_n169# 0 14.266f  
C475 a_864_n132# 0 30.763f  
C476 c3 0 23.08f  
C477 p3 0 0.378435p  
C478 a_579_n113# 0 18.082f  
C479 a_688_n102# 0 14.266f  
C480 a_302_n114# 0 30.763f  
C481 a_269_n114# 0 14.266f  
C482 a_324_n46# 0 26.066f  
C483 s2 0 3.76f  
C484 a_815_n46# 0 26.066f  
C485 b1 0 93.114f  
C486 a1 0 0.140495p  
C487 a_612_n65# 0 44.863f  
C488 a_924_n35# 0 14.266f  
C489 a_848_2# 0 30.763f  
C490 c2 0 23.08f  
C491 p2 0 0.505775p  
C492 a_582_25# 0 18.082f  
C493 a_691_36# 0 14.266f  
C494 a_302_20# 0 30.763f  
C495 a_269_20# 0 14.266f  
C496 a_324_88# 0 26.066f  
C497 b0 0 90.734f  
C498 a0 0 0.144276p  
C499 s1 0 3.76f  
C500 a_798_100# 0 26.066f  
C501 a_615_73# 0 44.863f  
C502 c1 0 23.08f  
C503 a_445_140# 0 4.888f  
C504 a_445_147# 0 20.28f  
C505 a_907_111# 0 14.266f  
C506 a_831_148# 0 30.763f  
C507 p1 0 0.380473p  
C508 pocin 0 28.03f  
C509 a_271_142# 0 18.082f  
C510 a_380_153# 0 14.266f  
C511 a_496_232# 0 1.316f  
C512 cin 0 85.827f  
C513 p0 0 0.200305p  
C514 s0 0 3.76f  
C515 a_738_234# 0 26.066f  
C516 a_304_190# 0 44.863f  
C517 a_496_251# 0 1.316f  
C518 p1p0c0 0 12.783999f  
C519 a_617_278# 0 4.888f  
C520 p1g0 0 18.06f  
C521 a_600_239# 0 21.819f  
C522 a_847_245# 0 14.266f  
C523 a_771_282# 0 30.763f  
C524 a_617_318# 0 2.585f  
C525 g1 0 0.241318p  
C526 a_453_311# 0 17.907999f  
C527 a_271_280# 0 18.082f  
C528 c4 0 4.324f  
C529 p3p2p1p0c0 0 12.783999f  
C530 a_380_291# 0 14.266f  
C531 a_610_377# 0 1.128f  
C532 g0 0 0.142494p  
C533 a_304_328# 0 44.863f  
C534 a_440_393# 0 1.316f  
C535 a_610_395# 0 1.316f  
C536 a_883_389# 0 4.888f  
C537 p3p2p1g0 0 18.624f  
C538 a_825_350# 0 23.605001f  
C539 p2g1 0 12.22f  
C540 a_610_414# 0 1.316f  
C541 a_440_412# 0 1.316f  
C542 a_731_417# 0 4.888f  
C543 p2p1p0c0 0 18.624f  
C544 a_883_429# 0 2.585f  
C545 p3p2g1 0 30.286f  
C546 a_693_378# 0 22.75f  
C547 a_731_457# 0 2.585f  
C548 p2p1g0 0 30.286f  
C549 a_883_464# 0 2.35f  
C550 p3g2 0 40.25f  
C551 a_218_418# 0 18.082f  
C552 a_534_474# 0 18.762999f  
C553 a_397_472# 0 17.907999f  
C554 a_327_429# 0 14.266f  
C555 a_731_492# 0 2.35f  
C556 g2 0 0.205115p  
C557 a_884_498# 0 2.115f  
C558 a_251_466# 0 44.863f  
C559 a_424_535# 0 1.316f  
C560 a_594_537# 0 1.316f  
C561 a_797_547# 0 1.316f  
C562 a_594_556# 0 1.316f  
C563 a_424_554# 0 1.316f  
C564 a_797_566# 0 1.316f  
C565 a_594_575# 0 1.316f  
C566 a_797_585# 0 1.316f  
C567 a_797_604# 0 1.316f  
C568 a_206_556# 0 18.082f  
C569 a_315_567# 0 14.266f  
C570 a_381_614# 0 17.907999f  
C571 a_239_604# 0 44.863f  
C572 a_518_635# 0 18.762999f  
C573 a_688_664# 0 19.618f  


 


* * RISING DELAY MEASUREMENT
* * Measure the delay for the final carry-out signal (C4)
.measure tran delay_C4 TRIG V(a0) VAL=0.9 RISE=1 TARG V(c4) VAL=0.9 RISE=1

* Measure the delay for each sum signal
.measure tran delay_S0 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s0) VAL=0.9 RISE=1
.measure tran delay_S1 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s1) VAL=0.9 RISE=1
.measure tran delay_S2 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s2) VAL=0.9 RISE=1
.measure tran delay_S3 TRIG V(a0) VAL=0.9 RISE=1 TARG V(s3) VAL=0.9 RISE=1


* FALLING DELAY MEASUREMENT
* Measure the delay for the final carry-out signal (C4)
* .measure tran delay_C4 TRIG V(a0) VAL=0.1 FALL=1 TARG V(c4) VAL=0.1 FALL=1

* * Measure the delay for each sum signal
* .measure tran delay_S0 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s0) VAL=0.1 FALL=1
* .measure tran delay_S1 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s1) VAL=0.1 FALL=1
* .measure tran delay_S2 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s2) VAL=0.1 FALL=1
* .measure tran delay_S3 TRIG V(a0) VAL=0.1 FALL=1 TARG V(s3) VAL=0.1 FALL=1




.control
  set hcopypscolor = 1             
  set color0 = white               
  set color1 = black               
  set color2 = red                 
  set color3 = blue                
  set color4 = coral               
  set color5 = brown    
  set color6 = cyan
  set color7 = chocolate   
  set color8 = chocolate
  set color9 = blueviolet
  set color10 = cadetblue        
  * for testing        
  * tran 1n 160n
  * for delay  
  tran 0.01n 20n 
   plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+g0 20+g1 22+g2 24+g3   
  plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+p0 20+p1 22+p2 24+p3                      
  plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+s0 20+s1 22+s2 24+s3                      
    plot a0 2+a1 4+a2 6+a3 8+b0 10+b1 12+b2 14+b3 16+cin 18+c4 20+s0 22+s1 24+s2 26+s3   
    * plot g3 2+p3g2 4+p3p2g1 6+p3p2p1g0 8+p3p2p1p0c0 10+c4 
    plot c1 2+p1 4+s1
  plot s0 2+s1 4+s2 6+s3    
        
.endc