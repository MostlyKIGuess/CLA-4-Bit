magic
tech scmos
timestamp 1731744794
<< nwell >>
rect 193 588 217 644
rect 226 594 250 650
rect 302 599 326 655
rect 335 599 359 655
rect 368 604 392 660
rect 401 604 425 660
rect 434 604 458 660
rect 472 604 496 660
rect 505 625 529 681
rect 538 625 562 681
rect 571 625 595 681
rect 604 625 628 681
rect 642 625 666 681
rect 675 654 699 710
rect 708 654 732 710
rect 741 654 765 710
rect 774 654 798 710
rect 807 654 831 710
rect 845 654 869 710
rect 205 450 229 506
rect 238 456 262 512
rect 314 461 338 517
rect 347 461 371 517
rect 384 462 408 518
rect 417 462 441 518
rect 450 462 474 518
rect 488 462 512 518
rect 521 464 545 520
rect 554 464 578 520
rect 587 464 611 520
rect 620 464 644 520
rect 658 464 682 520
rect 726 513 782 537
rect 879 518 935 542
rect 725 479 781 503
rect 878 485 934 509
rect 725 444 781 468
rect 725 411 781 435
rect 790 410 814 466
rect 877 451 933 475
rect 877 416 933 440
rect 877 383 933 407
rect 942 382 966 438
rect 258 312 282 368
rect 291 318 315 374
rect 367 323 391 379
rect 400 323 424 379
rect 440 301 464 357
rect 473 301 497 357
rect 506 301 530 357
rect 544 301 568 357
rect 611 340 667 364
rect 611 305 667 329
rect 611 272 667 296
rect 676 271 700 327
rect 725 266 749 322
rect 758 272 782 328
rect 797 280 821 332
rect 834 277 858 333
rect 867 277 891 333
rect 258 174 282 230
rect 291 180 315 236
rect 367 185 391 241
rect 400 185 424 241
rect 439 167 495 191
rect 439 134 495 158
rect 504 133 528 189
rect 258 17 282 73
rect 291 17 315 73
rect 328 18 352 70
rect 367 22 391 78
rect 400 28 424 84
rect 551 57 575 113
rect 584 63 608 119
rect 660 68 684 124
rect 693 68 717 124
rect 258 -117 282 -61
rect 291 -117 315 -61
rect 328 -116 352 -64
rect 367 -112 391 -56
rect 400 -106 424 -50
rect 548 -81 572 -25
rect 581 -75 605 -19
rect 657 -70 681 -14
rect 690 -70 714 -14
rect 785 -81 809 -25
rect 818 -75 842 -19
rect 857 -67 881 -15
rect 329 -250 353 -198
rect 368 -246 392 -190
rect 401 -240 425 -184
rect 551 -219 575 -163
rect 584 -213 608 -157
rect 782 -215 806 -159
rect 815 -209 839 -153
rect 854 -201 878 -149
rect 329 -384 353 -332
rect 368 -380 392 -324
rect 401 -374 425 -318
rect 551 -357 575 -301
rect 584 -351 608 -295
rect 660 -346 684 -290
rect 693 -346 717 -290
rect 795 -349 819 -293
rect 828 -343 852 -287
rect 867 -335 891 -283
<< ntransistor >>
rect 252 667 272 669
rect 797 621 837 623
rect 856 622 858 642
rect 252 581 272 583
rect 204 556 206 576
rect 313 567 315 587
rect 346 567 348 587
rect 424 571 464 573
rect 483 572 485 592
rect 594 592 634 594
rect 653 593 655 613
rect 797 602 837 604
rect 797 583 837 585
rect 594 573 634 575
rect 797 564 837 566
rect 424 552 464 554
rect 594 554 634 556
rect 797 545 837 547
rect 424 533 464 535
rect 594 535 634 537
rect 264 529 284 531
rect 264 443 284 445
rect 216 418 218 438
rect 325 429 327 449
rect 358 429 360 449
rect 440 429 480 431
rect 499 430 501 450
rect 610 431 650 433
rect 669 432 671 452
rect 440 410 480 412
rect 610 412 650 414
rect 317 391 337 393
rect 440 391 480 393
rect 610 393 650 395
rect 691 378 693 398
rect 712 378 714 398
rect 741 378 743 398
rect 774 378 776 398
rect 801 378 803 398
rect 610 375 650 377
rect 823 350 825 370
rect 843 350 845 370
rect 864 350 866 370
rect 893 350 895 370
rect 926 350 928 370
rect 953 350 955 370
rect 317 305 337 307
rect 269 280 271 300
rect 378 291 380 311
rect 411 291 413 311
rect 496 268 536 270
rect 555 269 557 289
rect 317 253 337 255
rect 496 249 536 251
rect 598 239 600 259
rect 627 239 629 259
rect 660 239 662 259
rect 687 239 689 259
rect 784 258 804 260
rect 736 234 738 254
rect 496 230 536 232
rect 821 233 823 253
rect 845 245 847 265
rect 878 245 880 265
rect 317 167 337 169
rect 269 142 271 162
rect 378 153 380 173
rect 411 153 413 173
rect 610 136 630 138
rect 269 85 271 105
rect 302 85 304 105
rect 326 97 328 117
rect 411 96 413 116
rect 455 101 457 121
rect 488 101 490 121
rect 515 101 517 121
rect 345 90 365 92
rect 610 50 630 52
rect 562 25 564 45
rect 671 36 673 56
rect 704 36 706 56
rect 607 -2 627 0
rect 269 -49 271 -29
rect 302 -49 304 -29
rect 326 -37 328 -17
rect 411 -38 413 -18
rect 345 -44 365 -42
rect 607 -88 627 -86
rect 559 -113 561 -93
rect 668 -102 670 -82
rect 701 -102 703 -82
rect 844 -89 864 -87
rect 796 -113 798 -93
rect 881 -114 883 -94
rect 610 -140 630 -138
rect 327 -171 329 -151
rect 412 -172 414 -152
rect 346 -178 366 -176
rect 610 -226 630 -224
rect 841 -223 861 -221
rect 562 -251 564 -231
rect 793 -247 795 -227
rect 878 -248 880 -228
rect 610 -278 630 -276
rect 327 -305 329 -285
rect 412 -306 414 -286
rect 346 -312 366 -310
rect 610 -364 630 -362
rect 562 -389 564 -369
rect 671 -378 673 -358
rect 704 -378 706 -358
rect 854 -357 874 -355
rect 806 -381 808 -361
rect 891 -382 893 -362
<< ptransistor >>
rect 204 598 206 638
rect 237 604 239 644
rect 313 609 315 649
rect 346 609 348 649
rect 379 614 381 654
rect 412 614 414 654
rect 445 614 447 654
rect 483 614 485 654
rect 516 635 518 675
rect 549 635 551 675
rect 582 635 584 675
rect 615 635 617 675
rect 653 635 655 675
rect 686 664 688 704
rect 719 664 721 704
rect 752 664 754 704
rect 785 664 787 704
rect 818 664 820 704
rect 856 664 858 704
rect 885 529 925 531
rect 732 524 772 526
rect 216 460 218 500
rect 249 466 251 506
rect 325 471 327 511
rect 358 471 360 511
rect 395 472 397 512
rect 428 472 430 512
rect 461 472 463 512
rect 499 472 501 512
rect 532 474 534 514
rect 565 474 567 514
rect 598 474 600 514
rect 631 474 633 514
rect 669 474 671 514
rect 884 496 924 498
rect 731 490 771 492
rect 883 462 923 464
rect 731 455 771 457
rect 731 422 771 424
rect 801 420 803 460
rect 883 427 923 429
rect 883 394 923 396
rect 953 392 955 432
rect 269 322 271 362
rect 302 328 304 368
rect 378 333 380 373
rect 411 333 413 373
rect 451 311 453 351
rect 484 311 486 351
rect 517 311 519 351
rect 555 311 557 351
rect 617 351 657 353
rect 617 316 657 318
rect 617 283 657 285
rect 687 281 689 321
rect 736 276 738 316
rect 769 282 771 322
rect 808 286 810 326
rect 845 287 847 327
rect 878 287 880 327
rect 269 184 271 224
rect 302 190 304 230
rect 378 195 380 235
rect 411 195 413 235
rect 445 178 485 180
rect 445 145 485 147
rect 515 143 517 183
rect 269 23 271 63
rect 302 23 304 63
rect 339 24 341 64
rect 378 28 380 68
rect 411 34 413 74
rect 562 67 564 107
rect 595 73 597 113
rect 671 78 673 118
rect 704 78 706 118
rect 269 -111 271 -71
rect 302 -111 304 -71
rect 339 -110 341 -70
rect 378 -106 380 -66
rect 411 -100 413 -60
rect 559 -71 561 -31
rect 592 -65 594 -25
rect 668 -60 670 -20
rect 701 -60 703 -20
rect 796 -71 798 -31
rect 829 -65 831 -25
rect 868 -61 870 -21
rect 340 -244 342 -204
rect 379 -240 381 -200
rect 412 -234 414 -194
rect 562 -209 564 -169
rect 595 -203 597 -163
rect 793 -205 795 -165
rect 826 -199 828 -159
rect 865 -195 867 -155
rect 340 -378 342 -338
rect 379 -374 381 -334
rect 412 -368 414 -328
rect 562 -347 564 -307
rect 595 -341 597 -301
rect 671 -336 673 -296
rect 704 -336 706 -296
rect 806 -339 808 -299
rect 839 -333 841 -293
rect 878 -329 880 -289
<< ndiffusion >>
rect 252 669 272 670
rect 252 666 272 667
rect 797 623 837 624
rect 855 622 856 642
rect 858 622 859 642
rect 797 620 837 621
rect 252 583 272 584
rect 252 580 272 581
rect 203 556 204 576
rect 206 556 207 576
rect 312 567 313 587
rect 315 567 316 587
rect 345 567 346 587
rect 348 567 349 587
rect 424 573 464 574
rect 482 572 483 592
rect 485 572 486 592
rect 594 594 634 595
rect 652 593 653 613
rect 655 593 656 613
rect 797 604 837 605
rect 797 601 837 602
rect 594 591 634 592
rect 797 585 837 586
rect 797 582 837 583
rect 424 570 464 571
rect 594 575 634 576
rect 594 572 634 573
rect 797 566 837 567
rect 797 563 837 564
rect 424 554 464 555
rect 594 556 634 557
rect 594 553 634 554
rect 424 551 464 552
rect 797 547 837 548
rect 797 544 837 545
rect 264 531 284 532
rect 424 535 464 536
rect 594 537 634 538
rect 594 534 634 535
rect 424 532 464 533
rect 264 528 284 529
rect 264 445 284 446
rect 264 442 284 443
rect 215 418 216 438
rect 218 418 219 438
rect 324 429 325 449
rect 327 429 328 449
rect 357 429 358 449
rect 360 429 361 449
rect 440 431 480 432
rect 498 430 499 450
rect 501 430 502 450
rect 440 428 480 429
rect 610 433 650 434
rect 668 432 669 452
rect 671 432 672 452
rect 610 430 650 431
rect 440 412 480 413
rect 610 414 650 415
rect 610 411 650 412
rect 440 409 480 410
rect 317 393 337 394
rect 317 390 337 391
rect 440 393 480 394
rect 610 395 650 396
rect 610 392 650 393
rect 440 390 480 391
rect 690 378 691 398
rect 693 378 694 398
rect 711 378 712 398
rect 714 378 715 398
rect 740 378 741 398
rect 743 378 744 398
rect 773 378 774 398
rect 776 378 777 398
rect 800 378 801 398
rect 803 378 804 398
rect 610 377 650 378
rect 610 374 650 375
rect 822 350 823 370
rect 825 350 826 370
rect 842 350 843 370
rect 845 350 846 370
rect 863 350 864 370
rect 866 350 867 370
rect 892 350 893 370
rect 895 350 896 370
rect 925 350 926 370
rect 928 350 929 370
rect 952 350 953 370
rect 955 350 956 370
rect 317 307 337 308
rect 317 304 337 305
rect 268 280 269 300
rect 271 280 272 300
rect 377 291 378 311
rect 380 291 381 311
rect 410 291 411 311
rect 413 291 414 311
rect 496 270 536 271
rect 554 269 555 289
rect 557 269 558 289
rect 496 267 536 268
rect 317 255 337 256
rect 317 252 337 253
rect 496 251 536 252
rect 496 248 536 249
rect 597 239 598 259
rect 600 239 601 259
rect 626 239 627 259
rect 629 239 630 259
rect 659 239 660 259
rect 662 239 663 259
rect 686 239 687 259
rect 689 239 690 259
rect 784 260 804 261
rect 784 257 804 258
rect 735 234 736 254
rect 738 234 739 254
rect 496 232 536 233
rect 820 233 821 253
rect 823 233 824 253
rect 844 245 845 265
rect 847 245 848 265
rect 877 245 878 265
rect 880 245 881 265
rect 496 229 536 230
rect 317 169 337 170
rect 317 166 337 167
rect 268 142 269 162
rect 271 142 272 162
rect 377 153 378 173
rect 380 153 381 173
rect 410 153 411 173
rect 413 153 414 173
rect 610 138 630 139
rect 610 135 630 136
rect 268 85 269 105
rect 271 85 272 105
rect 301 85 302 105
rect 304 85 305 105
rect 325 97 326 117
rect 328 97 329 117
rect 410 96 411 116
rect 413 96 414 116
rect 454 101 455 121
rect 457 101 458 121
rect 487 101 488 121
rect 490 101 491 121
rect 514 101 515 121
rect 517 101 518 121
rect 345 92 365 93
rect 345 89 365 90
rect 610 52 630 53
rect 610 49 630 50
rect 561 25 562 45
rect 564 25 565 45
rect 670 36 671 56
rect 673 36 674 56
rect 703 36 704 56
rect 706 36 707 56
rect 607 0 627 1
rect 607 -3 627 -2
rect 268 -49 269 -29
rect 271 -49 272 -29
rect 301 -49 302 -29
rect 304 -49 305 -29
rect 325 -37 326 -17
rect 328 -37 329 -17
rect 410 -38 411 -18
rect 413 -38 414 -18
rect 345 -42 365 -41
rect 345 -45 365 -44
rect 607 -86 627 -85
rect 607 -89 627 -88
rect 558 -113 559 -93
rect 561 -113 562 -93
rect 667 -102 668 -82
rect 670 -102 671 -82
rect 700 -102 701 -82
rect 703 -102 704 -82
rect 844 -87 864 -86
rect 844 -90 864 -89
rect 795 -113 796 -93
rect 798 -113 799 -93
rect 880 -114 881 -94
rect 883 -114 884 -94
rect 610 -138 630 -137
rect 610 -141 630 -140
rect 326 -171 327 -151
rect 329 -171 330 -151
rect 411 -172 412 -152
rect 414 -172 415 -152
rect 346 -176 366 -175
rect 346 -179 366 -178
rect 610 -224 630 -223
rect 610 -227 630 -226
rect 841 -221 861 -220
rect 841 -224 861 -223
rect 561 -251 562 -231
rect 564 -251 565 -231
rect 792 -247 793 -227
rect 795 -247 796 -227
rect 877 -248 878 -228
rect 880 -248 881 -228
rect 610 -276 630 -275
rect 610 -279 630 -278
rect 326 -305 327 -285
rect 329 -305 330 -285
rect 411 -306 412 -286
rect 414 -306 415 -286
rect 346 -310 366 -309
rect 346 -313 366 -312
rect 610 -362 630 -361
rect 610 -365 630 -364
rect 561 -389 562 -369
rect 564 -389 565 -369
rect 670 -378 671 -358
rect 673 -378 674 -358
rect 703 -378 704 -358
rect 706 -378 707 -358
rect 854 -355 874 -354
rect 854 -358 874 -357
rect 805 -381 806 -361
rect 808 -381 809 -361
rect 890 -382 891 -362
rect 893 -382 894 -362
<< pdiffusion >>
rect 203 598 204 638
rect 206 598 207 638
rect 236 604 237 644
rect 239 604 240 644
rect 312 609 313 649
rect 315 609 316 649
rect 345 609 346 649
rect 348 609 349 649
rect 378 614 379 654
rect 381 614 382 654
rect 411 614 412 654
rect 414 614 415 654
rect 444 614 445 654
rect 447 614 448 654
rect 482 614 483 654
rect 485 614 486 654
rect 515 635 516 675
rect 518 635 519 675
rect 548 635 549 675
rect 551 635 552 675
rect 581 635 582 675
rect 584 635 585 675
rect 614 635 615 675
rect 617 635 618 675
rect 652 635 653 675
rect 655 635 656 675
rect 685 664 686 704
rect 688 664 689 704
rect 718 664 719 704
rect 721 664 722 704
rect 751 664 752 704
rect 754 664 755 704
rect 784 664 785 704
rect 787 664 788 704
rect 817 664 818 704
rect 820 664 821 704
rect 855 664 856 704
rect 858 664 859 704
rect 885 531 925 532
rect 885 528 925 529
rect 732 526 772 527
rect 732 523 772 524
rect 215 460 216 500
rect 218 460 219 500
rect 248 466 249 506
rect 251 466 252 506
rect 324 471 325 511
rect 327 471 328 511
rect 357 471 358 511
rect 360 471 361 511
rect 394 472 395 512
rect 397 472 398 512
rect 427 472 428 512
rect 430 472 431 512
rect 460 472 461 512
rect 463 472 464 512
rect 498 472 499 512
rect 501 472 502 512
rect 531 474 532 514
rect 534 474 535 514
rect 564 474 565 514
rect 567 474 568 514
rect 597 474 598 514
rect 600 474 601 514
rect 630 474 631 514
rect 633 474 634 514
rect 668 474 669 514
rect 671 474 672 514
rect 884 498 924 499
rect 884 495 924 496
rect 731 492 771 493
rect 731 489 771 490
rect 883 464 923 465
rect 883 461 923 462
rect 731 457 771 458
rect 731 454 771 455
rect 731 424 771 425
rect 731 421 771 422
rect 800 420 801 460
rect 803 420 804 460
rect 883 429 923 430
rect 883 426 923 427
rect 883 396 923 397
rect 883 393 923 394
rect 952 392 953 432
rect 955 392 956 432
rect 268 322 269 362
rect 271 322 272 362
rect 301 328 302 368
rect 304 328 305 368
rect 377 333 378 373
rect 380 333 381 373
rect 410 333 411 373
rect 413 333 414 373
rect 450 311 451 351
rect 453 311 454 351
rect 483 311 484 351
rect 486 311 487 351
rect 516 311 517 351
rect 519 311 520 351
rect 554 311 555 351
rect 557 311 558 351
rect 617 353 657 354
rect 617 350 657 351
rect 617 318 657 319
rect 617 315 657 316
rect 617 285 657 286
rect 617 282 657 283
rect 686 281 687 321
rect 689 281 690 321
rect 735 276 736 316
rect 738 276 739 316
rect 768 282 769 322
rect 771 282 772 322
rect 807 286 808 326
rect 810 286 811 326
rect 844 287 845 327
rect 847 287 848 327
rect 877 287 878 327
rect 880 287 881 327
rect 268 184 269 224
rect 271 184 272 224
rect 301 190 302 230
rect 304 190 305 230
rect 377 195 378 235
rect 380 195 381 235
rect 410 195 411 235
rect 413 195 414 235
rect 445 180 485 181
rect 445 177 485 178
rect 445 147 485 148
rect 445 144 485 145
rect 514 143 515 183
rect 517 143 518 183
rect 268 23 269 63
rect 271 23 272 63
rect 301 23 302 63
rect 304 23 305 63
rect 338 24 339 64
rect 341 24 342 64
rect 377 28 378 68
rect 380 28 381 68
rect 410 34 411 74
rect 413 34 414 74
rect 561 67 562 107
rect 564 67 565 107
rect 594 73 595 113
rect 597 73 598 113
rect 670 78 671 118
rect 673 78 674 118
rect 703 78 704 118
rect 706 78 707 118
rect 268 -111 269 -71
rect 271 -111 272 -71
rect 301 -111 302 -71
rect 304 -111 305 -71
rect 338 -110 339 -70
rect 341 -110 342 -70
rect 377 -106 378 -66
rect 380 -106 381 -66
rect 410 -100 411 -60
rect 413 -100 414 -60
rect 558 -71 559 -31
rect 561 -71 562 -31
rect 591 -65 592 -25
rect 594 -65 595 -25
rect 667 -60 668 -20
rect 670 -60 671 -20
rect 700 -60 701 -20
rect 703 -60 704 -20
rect 795 -71 796 -31
rect 798 -71 799 -31
rect 828 -65 829 -25
rect 831 -65 832 -25
rect 867 -61 868 -21
rect 870 -61 871 -21
rect 339 -244 340 -204
rect 342 -244 343 -204
rect 378 -240 379 -200
rect 381 -240 382 -200
rect 411 -234 412 -194
rect 414 -234 415 -194
rect 561 -209 562 -169
rect 564 -209 565 -169
rect 594 -203 595 -163
rect 597 -203 598 -163
rect 792 -205 793 -165
rect 795 -205 796 -165
rect 825 -199 826 -159
rect 828 -199 829 -159
rect 864 -195 865 -155
rect 867 -195 868 -155
rect 339 -378 340 -338
rect 342 -378 343 -338
rect 378 -374 379 -334
rect 381 -374 382 -334
rect 411 -368 412 -328
rect 414 -368 415 -328
rect 561 -347 562 -307
rect 564 -347 565 -307
rect 594 -341 595 -301
rect 597 -341 598 -301
rect 670 -336 671 -296
rect 673 -336 674 -296
rect 703 -336 704 -296
rect 706 -336 707 -296
rect 805 -339 806 -299
rect 808 -339 809 -299
rect 838 -333 839 -293
rect 841 -333 842 -293
rect 877 -329 878 -289
rect 880 -329 881 -289
<< ndcontact >>
rect 252 670 272 674
rect 252 662 272 666
rect 252 584 272 588
rect 797 624 837 628
rect 851 622 855 642
rect 859 622 863 642
rect 797 616 837 620
rect 252 576 272 580
rect 199 556 203 576
rect 207 556 211 576
rect 308 567 312 587
rect 316 567 320 587
rect 341 567 345 587
rect 349 567 353 587
rect 424 574 464 578
rect 478 572 482 592
rect 486 572 490 592
rect 594 595 634 599
rect 648 593 652 613
rect 656 593 660 613
rect 797 605 837 609
rect 797 597 837 601
rect 594 587 634 591
rect 797 586 837 590
rect 424 566 464 570
rect 594 576 634 580
rect 797 578 837 582
rect 594 568 634 572
rect 797 567 837 571
rect 424 555 464 559
rect 594 557 634 561
rect 797 559 837 563
rect 424 547 464 551
rect 594 549 634 553
rect 797 548 837 552
rect 264 532 284 536
rect 424 536 464 540
rect 594 538 634 542
rect 797 540 837 544
rect 424 528 464 532
rect 594 530 634 534
rect 264 524 284 528
rect 264 446 284 450
rect 264 438 284 442
rect 211 418 215 438
rect 219 418 223 438
rect 320 429 324 449
rect 328 429 332 449
rect 353 429 357 449
rect 361 429 365 449
rect 440 432 480 436
rect 494 430 498 450
rect 502 430 506 450
rect 440 424 480 428
rect 610 434 650 438
rect 664 432 668 452
rect 672 432 676 452
rect 610 426 650 430
rect 440 413 480 417
rect 610 415 650 419
rect 440 405 480 409
rect 610 407 650 411
rect 317 394 337 398
rect 317 386 337 390
rect 440 394 480 398
rect 610 396 650 400
rect 440 386 480 390
rect 610 388 650 392
rect 610 378 650 382
rect 686 378 690 398
rect 694 378 698 398
rect 707 378 711 398
rect 715 378 719 398
rect 736 378 740 398
rect 744 378 748 398
rect 769 378 773 398
rect 777 378 781 398
rect 796 378 800 398
rect 804 378 808 398
rect 610 370 650 374
rect 317 308 337 312
rect 818 350 822 370
rect 826 350 830 370
rect 838 350 842 370
rect 846 350 850 370
rect 859 350 863 370
rect 867 350 871 370
rect 888 350 892 370
rect 896 350 900 370
rect 921 350 925 370
rect 929 350 933 370
rect 948 350 952 370
rect 956 350 960 370
rect 317 300 337 304
rect 264 280 268 300
rect 272 280 276 300
rect 373 291 377 311
rect 381 291 385 311
rect 406 291 410 311
rect 414 291 418 311
rect 496 271 536 275
rect 550 269 554 289
rect 558 269 562 289
rect 496 263 536 267
rect 317 256 337 260
rect 317 248 337 252
rect 496 252 536 256
rect 496 244 536 248
rect 593 239 597 259
rect 601 239 605 259
rect 622 239 626 259
rect 630 239 634 259
rect 655 239 659 259
rect 663 239 667 259
rect 682 239 686 259
rect 690 239 694 259
rect 784 261 804 265
rect 496 233 536 237
rect 731 234 735 254
rect 739 234 743 254
rect 784 253 804 257
rect 816 233 820 253
rect 824 233 828 253
rect 840 245 844 265
rect 848 245 852 265
rect 873 245 877 265
rect 881 245 885 265
rect 496 225 536 229
rect 317 170 337 174
rect 317 162 337 166
rect 264 142 268 162
rect 272 142 276 162
rect 373 153 377 173
rect 381 153 385 173
rect 406 153 410 173
rect 414 153 418 173
rect 610 139 630 143
rect 610 131 630 135
rect 264 85 268 105
rect 272 85 276 105
rect 297 85 301 105
rect 305 85 309 105
rect 321 97 325 117
rect 329 97 333 117
rect 345 93 365 97
rect 406 96 410 116
rect 414 96 418 116
rect 450 101 454 121
rect 458 101 462 121
rect 483 101 487 121
rect 491 101 495 121
rect 510 101 514 121
rect 518 101 522 121
rect 345 85 365 89
rect 610 53 630 57
rect 610 45 630 49
rect 557 25 561 45
rect 565 25 569 45
rect 666 36 670 56
rect 674 36 678 56
rect 699 36 703 56
rect 707 36 711 56
rect 607 1 627 5
rect 607 -7 627 -3
rect 264 -49 268 -29
rect 272 -49 276 -29
rect 297 -49 301 -29
rect 305 -49 309 -29
rect 321 -37 325 -17
rect 329 -37 333 -17
rect 345 -41 365 -37
rect 406 -38 410 -18
rect 414 -38 418 -18
rect 345 -49 365 -45
rect 607 -85 627 -81
rect 607 -93 627 -89
rect 554 -113 558 -93
rect 562 -113 566 -93
rect 663 -102 667 -82
rect 671 -102 675 -82
rect 696 -102 700 -82
rect 704 -102 708 -82
rect 844 -86 864 -82
rect 791 -113 795 -93
rect 799 -113 803 -93
rect 844 -94 864 -90
rect 876 -114 880 -94
rect 884 -114 888 -94
rect 610 -137 630 -133
rect 610 -145 630 -141
rect 322 -171 326 -151
rect 330 -171 334 -151
rect 346 -175 366 -171
rect 407 -172 411 -152
rect 415 -172 419 -152
rect 346 -183 366 -179
rect 610 -223 630 -219
rect 841 -220 861 -216
rect 610 -231 630 -227
rect 557 -251 561 -231
rect 565 -251 569 -231
rect 788 -247 792 -227
rect 796 -247 800 -227
rect 841 -228 861 -224
rect 873 -248 877 -228
rect 881 -248 885 -228
rect 610 -275 630 -271
rect 610 -283 630 -279
rect 322 -305 326 -285
rect 330 -305 334 -285
rect 346 -309 366 -305
rect 407 -306 411 -286
rect 415 -306 419 -286
rect 346 -317 366 -313
rect 610 -361 630 -357
rect 610 -369 630 -365
rect 557 -389 561 -369
rect 565 -389 569 -369
rect 666 -378 670 -358
rect 674 -378 678 -358
rect 699 -378 703 -358
rect 707 -378 711 -358
rect 854 -354 874 -350
rect 801 -381 805 -361
rect 809 -381 813 -361
rect 854 -362 874 -358
rect 886 -382 890 -362
rect 894 -382 898 -362
<< pdcontact >>
rect 199 598 203 638
rect 207 598 211 638
rect 232 604 236 644
rect 240 604 244 644
rect 308 609 312 649
rect 316 609 320 649
rect 341 609 345 649
rect 349 609 353 649
rect 374 614 378 654
rect 382 614 386 654
rect 407 614 411 654
rect 415 614 419 654
rect 440 614 444 654
rect 448 614 452 654
rect 478 614 482 654
rect 486 614 490 654
rect 511 635 515 675
rect 519 635 523 675
rect 544 635 548 675
rect 552 635 556 675
rect 577 635 581 675
rect 585 635 589 675
rect 610 635 614 675
rect 618 635 622 675
rect 648 635 652 675
rect 656 635 660 675
rect 681 664 685 704
rect 689 664 693 704
rect 714 664 718 704
rect 722 664 726 704
rect 747 664 751 704
rect 755 664 759 704
rect 780 664 784 704
rect 788 664 792 704
rect 813 664 817 704
rect 821 664 825 704
rect 851 664 855 704
rect 859 664 863 704
rect 885 532 925 536
rect 732 527 772 531
rect 885 524 925 528
rect 732 519 772 523
rect 211 460 215 500
rect 219 460 223 500
rect 244 466 248 506
rect 252 466 256 506
rect 320 471 324 511
rect 328 471 332 511
rect 353 471 357 511
rect 361 471 365 511
rect 390 472 394 512
rect 398 472 402 512
rect 423 472 427 512
rect 431 472 435 512
rect 456 472 460 512
rect 464 472 468 512
rect 494 472 498 512
rect 502 472 506 512
rect 527 474 531 514
rect 535 474 539 514
rect 560 474 564 514
rect 568 474 572 514
rect 593 474 597 514
rect 601 474 605 514
rect 626 474 630 514
rect 634 474 638 514
rect 664 474 668 514
rect 672 474 676 514
rect 884 499 924 503
rect 731 493 771 497
rect 884 491 924 495
rect 731 485 771 489
rect 883 465 923 469
rect 731 458 771 462
rect 731 450 771 454
rect 731 425 771 429
rect 731 417 771 421
rect 796 420 800 460
rect 804 420 808 460
rect 883 457 923 461
rect 883 430 923 434
rect 883 422 923 426
rect 883 397 923 401
rect 883 389 923 393
rect 948 392 952 432
rect 956 392 960 432
rect 264 322 268 362
rect 272 322 276 362
rect 297 328 301 368
rect 305 328 309 368
rect 373 333 377 373
rect 381 333 385 373
rect 406 333 410 373
rect 414 333 418 373
rect 617 354 657 358
rect 446 311 450 351
rect 454 311 458 351
rect 479 311 483 351
rect 487 311 491 351
rect 512 311 516 351
rect 520 311 524 351
rect 550 311 554 351
rect 558 311 562 351
rect 617 346 657 350
rect 617 319 657 323
rect 617 311 657 315
rect 617 286 657 290
rect 617 278 657 282
rect 682 281 686 321
rect 690 281 694 321
rect 731 276 735 316
rect 739 276 743 316
rect 764 282 768 322
rect 772 282 776 322
rect 803 286 807 326
rect 811 286 815 326
rect 840 287 844 327
rect 848 287 852 327
rect 873 287 877 327
rect 881 287 885 327
rect 264 184 268 224
rect 272 184 276 224
rect 297 190 301 230
rect 305 190 309 230
rect 373 195 377 235
rect 381 195 385 235
rect 406 195 410 235
rect 414 195 418 235
rect 445 181 485 185
rect 445 173 485 177
rect 445 148 485 152
rect 445 140 485 144
rect 510 143 514 183
rect 518 143 522 183
rect 264 23 268 63
rect 272 23 276 63
rect 297 23 301 63
rect 305 23 309 63
rect 334 24 338 64
rect 342 24 346 64
rect 373 28 377 68
rect 381 28 385 68
rect 406 34 410 74
rect 414 34 418 74
rect 557 67 561 107
rect 565 67 569 107
rect 590 73 594 113
rect 598 73 602 113
rect 666 78 670 118
rect 674 78 678 118
rect 699 78 703 118
rect 707 78 711 118
rect 264 -111 268 -71
rect 272 -111 276 -71
rect 297 -111 301 -71
rect 305 -111 309 -71
rect 334 -110 338 -70
rect 342 -110 346 -70
rect 373 -106 377 -66
rect 381 -106 385 -66
rect 406 -100 410 -60
rect 414 -100 418 -60
rect 554 -71 558 -31
rect 562 -71 566 -31
rect 587 -65 591 -25
rect 595 -65 599 -25
rect 663 -60 667 -20
rect 671 -60 675 -20
rect 696 -60 700 -20
rect 704 -60 708 -20
rect 791 -71 795 -31
rect 799 -71 803 -31
rect 824 -65 828 -25
rect 832 -65 836 -25
rect 863 -61 867 -21
rect 871 -61 875 -21
rect 335 -244 339 -204
rect 343 -244 347 -204
rect 374 -240 378 -200
rect 382 -240 386 -200
rect 407 -234 411 -194
rect 415 -234 419 -194
rect 557 -209 561 -169
rect 565 -209 569 -169
rect 590 -203 594 -163
rect 598 -203 602 -163
rect 788 -205 792 -165
rect 796 -205 800 -165
rect 821 -199 825 -159
rect 829 -199 833 -159
rect 860 -195 864 -155
rect 868 -195 872 -155
rect 335 -378 339 -338
rect 343 -378 347 -338
rect 374 -374 378 -334
rect 382 -374 386 -334
rect 407 -368 411 -328
rect 415 -368 419 -328
rect 557 -347 561 -307
rect 565 -347 569 -307
rect 590 -341 594 -301
rect 598 -341 602 -301
rect 666 -336 670 -296
rect 674 -336 678 -296
rect 699 -336 703 -296
rect 707 -336 711 -296
rect 801 -339 805 -299
rect 809 -339 813 -299
rect 834 -333 838 -293
rect 842 -333 846 -293
rect 873 -329 877 -289
rect 881 -329 885 -289
<< polysilicon >>
rect 686 704 688 707
rect 719 704 721 707
rect 752 704 754 707
rect 785 704 787 707
rect 818 704 820 707
rect 856 704 858 707
rect 516 675 518 678
rect 549 675 551 678
rect 582 675 584 678
rect 615 675 617 678
rect 653 675 655 678
rect 249 667 252 669
rect 272 667 275 669
rect 379 654 381 657
rect 412 654 414 657
rect 445 654 447 657
rect 483 654 485 657
rect 313 649 315 652
rect 346 649 348 652
rect 237 644 239 647
rect 204 638 206 641
rect 686 651 688 664
rect 719 651 721 664
rect 752 651 754 664
rect 785 651 787 664
rect 818 651 820 664
rect 856 642 858 664
rect 516 622 518 635
rect 549 622 551 635
rect 582 622 584 635
rect 615 622 617 635
rect 204 576 206 598
rect 237 592 239 604
rect 313 587 315 609
rect 346 587 348 609
rect 379 601 381 614
rect 412 601 414 614
rect 445 601 447 614
rect 483 592 485 614
rect 653 613 655 635
rect 794 621 797 623
rect 837 621 840 623
rect 856 619 858 622
rect 244 581 252 583
rect 272 581 275 583
rect 421 571 424 573
rect 464 571 467 573
rect 591 592 594 594
rect 634 592 637 594
rect 794 602 797 604
rect 837 602 840 604
rect 653 590 655 593
rect 794 583 797 585
rect 837 583 840 585
rect 313 564 315 567
rect 346 564 348 567
rect 483 569 485 572
rect 591 573 594 575
rect 634 573 637 575
rect 794 564 797 566
rect 837 564 840 566
rect 204 553 206 556
rect 421 552 424 554
rect 464 552 467 554
rect 591 554 594 556
rect 634 554 637 556
rect 794 545 797 547
rect 837 545 840 547
rect 421 533 424 535
rect 464 533 467 535
rect 591 535 594 537
rect 634 535 637 537
rect 261 529 264 531
rect 284 529 287 531
rect 882 529 885 531
rect 925 529 936 531
rect 729 524 732 526
rect 772 524 783 526
rect 325 511 327 514
rect 358 511 360 514
rect 395 512 397 515
rect 428 512 430 515
rect 461 512 463 515
rect 499 512 501 515
rect 532 514 534 517
rect 565 514 567 517
rect 598 514 600 517
rect 631 514 633 517
rect 669 514 671 517
rect 249 506 251 509
rect 216 500 218 503
rect 881 496 884 498
rect 924 496 935 498
rect 728 490 731 492
rect 771 490 782 492
rect 216 438 218 460
rect 249 454 251 466
rect 325 449 327 471
rect 358 449 360 471
rect 395 459 397 472
rect 428 459 430 472
rect 461 459 463 472
rect 499 450 501 472
rect 532 461 534 474
rect 565 461 567 474
rect 598 461 600 474
rect 631 461 633 474
rect 669 452 671 474
rect 801 460 803 463
rect 880 462 883 464
rect 923 462 934 464
rect 728 455 731 457
rect 771 455 782 457
rect 256 443 264 445
rect 284 443 287 445
rect 325 426 327 429
rect 358 426 360 429
rect 437 429 440 431
rect 480 429 483 431
rect 499 427 501 430
rect 607 431 610 433
rect 650 431 653 433
rect 669 429 671 432
rect 728 422 731 424
rect 771 422 777 424
rect 216 415 218 418
rect 437 410 440 412
rect 480 410 483 412
rect 775 418 777 422
rect 953 432 955 435
rect 880 427 883 429
rect 923 427 934 429
rect 607 412 610 414
rect 650 412 653 414
rect 314 391 317 393
rect 337 391 340 393
rect 437 391 440 393
rect 480 391 483 393
rect 691 398 693 401
rect 712 398 714 401
rect 741 398 743 401
rect 774 398 776 401
rect 801 398 803 420
rect 607 393 610 395
rect 650 393 653 395
rect 378 373 380 376
rect 411 373 413 376
rect 880 394 883 396
rect 923 394 929 396
rect 927 390 929 394
rect 607 375 610 377
rect 650 375 653 377
rect 691 375 693 378
rect 712 375 714 378
rect 741 375 743 378
rect 774 375 776 378
rect 801 375 803 378
rect 302 368 304 371
rect 269 362 271 365
rect 823 370 825 373
rect 843 370 845 373
rect 864 370 866 373
rect 893 370 895 373
rect 926 370 928 373
rect 953 370 955 392
rect 451 351 453 354
rect 484 351 486 354
rect 517 351 519 354
rect 555 351 557 354
rect 269 300 271 322
rect 302 316 304 328
rect 378 311 380 333
rect 411 311 413 333
rect 614 351 617 353
rect 657 351 668 353
rect 823 347 825 350
rect 843 347 845 350
rect 864 347 866 350
rect 893 347 895 350
rect 926 347 928 350
rect 953 347 955 350
rect 808 326 810 329
rect 845 327 847 330
rect 878 327 880 330
rect 687 321 689 324
rect 769 322 771 325
rect 614 316 617 318
rect 657 316 668 318
rect 309 305 317 307
rect 337 305 340 307
rect 451 298 453 311
rect 484 298 486 311
rect 517 298 519 311
rect 378 288 380 291
rect 411 288 413 291
rect 555 289 557 311
rect 269 277 271 280
rect 493 268 496 270
rect 536 268 539 270
rect 614 283 617 285
rect 657 283 663 285
rect 661 279 663 283
rect 736 316 738 319
rect 555 266 557 269
rect 598 259 600 262
rect 627 259 629 262
rect 660 259 662 262
rect 687 259 689 281
rect 808 283 810 286
rect 769 276 771 282
rect 314 253 317 255
rect 337 253 340 255
rect 493 249 496 251
rect 536 249 539 251
rect 736 254 738 276
rect 845 265 847 287
rect 878 265 880 287
rect 776 258 784 260
rect 804 258 807 260
rect 378 235 380 238
rect 411 235 413 238
rect 302 230 304 233
rect 269 224 271 227
rect 598 236 600 239
rect 627 236 629 239
rect 660 236 662 239
rect 687 236 689 239
rect 821 253 823 257
rect 493 230 496 232
rect 536 230 539 232
rect 736 231 738 234
rect 845 242 847 245
rect 878 242 880 245
rect 821 230 823 233
rect 269 162 271 184
rect 302 178 304 190
rect 378 173 380 195
rect 411 173 413 195
rect 515 183 517 186
rect 442 178 445 180
rect 485 178 496 180
rect 309 167 317 169
rect 337 167 340 169
rect 378 150 380 153
rect 411 150 413 153
rect 442 145 445 147
rect 485 145 491 147
rect 269 139 271 142
rect 489 141 491 145
rect 455 121 457 124
rect 488 121 490 124
rect 515 121 517 143
rect 607 136 610 138
rect 630 136 633 138
rect 326 117 328 120
rect 269 105 271 108
rect 302 105 304 108
rect 411 116 413 119
rect 326 93 328 97
rect 671 118 673 121
rect 704 118 706 121
rect 595 113 597 116
rect 562 107 564 110
rect 455 98 457 101
rect 488 98 490 101
rect 515 98 517 101
rect 342 90 345 92
rect 365 90 373 92
rect 269 63 271 85
rect 302 63 304 85
rect 411 74 413 96
rect 378 68 380 74
rect 339 64 341 67
rect 562 45 564 67
rect 595 61 597 73
rect 671 56 673 78
rect 704 56 706 78
rect 602 50 610 52
rect 630 50 633 52
rect 411 31 413 34
rect 378 25 380 28
rect 671 33 673 36
rect 704 33 706 36
rect 269 20 271 23
rect 302 20 304 23
rect 339 21 341 24
rect 562 22 564 25
rect 604 -2 607 0
rect 627 -2 630 0
rect 326 -17 328 -14
rect 269 -29 271 -26
rect 302 -29 304 -26
rect 411 -18 413 -15
rect 326 -41 328 -37
rect 668 -20 670 -17
rect 701 -20 703 -17
rect 592 -25 594 -22
rect 559 -31 561 -28
rect 342 -44 345 -42
rect 365 -44 373 -42
rect 269 -71 271 -49
rect 302 -71 304 -49
rect 411 -60 413 -38
rect 378 -66 380 -60
rect 339 -70 341 -67
rect 868 -21 870 -18
rect 829 -25 831 -22
rect 796 -31 798 -28
rect 559 -93 561 -71
rect 592 -77 594 -65
rect 668 -82 670 -60
rect 701 -82 703 -60
rect 868 -64 870 -61
rect 829 -71 831 -65
rect 599 -88 607 -86
rect 627 -88 630 -86
rect 411 -103 413 -100
rect 378 -109 380 -106
rect 269 -114 271 -111
rect 302 -114 304 -111
rect 339 -113 341 -110
rect 796 -93 798 -71
rect 836 -89 844 -87
rect 864 -89 867 -87
rect 668 -105 670 -102
rect 701 -105 703 -102
rect 881 -94 883 -90
rect 559 -116 561 -113
rect 796 -116 798 -113
rect 881 -117 883 -114
rect 607 -140 610 -138
rect 630 -140 633 -138
rect 327 -151 329 -148
rect 412 -152 414 -149
rect 327 -175 329 -171
rect 865 -155 867 -152
rect 826 -159 828 -156
rect 595 -163 597 -160
rect 562 -169 564 -166
rect 343 -178 346 -176
rect 366 -178 374 -176
rect 412 -194 414 -172
rect 379 -200 381 -194
rect 340 -204 342 -201
rect 793 -165 795 -162
rect 562 -231 564 -209
rect 595 -215 597 -203
rect 865 -198 867 -195
rect 826 -205 828 -199
rect 602 -226 610 -224
rect 630 -226 633 -224
rect 793 -227 795 -205
rect 833 -223 841 -221
rect 861 -223 864 -221
rect 412 -237 414 -234
rect 379 -243 381 -240
rect 340 -247 342 -244
rect 878 -228 880 -224
rect 793 -250 795 -247
rect 878 -251 880 -248
rect 562 -254 564 -251
rect 607 -278 610 -276
rect 630 -278 633 -276
rect 327 -285 329 -282
rect 412 -286 414 -283
rect 327 -309 329 -305
rect 878 -289 880 -286
rect 839 -293 841 -290
rect 671 -296 673 -293
rect 704 -296 706 -293
rect 595 -301 597 -298
rect 343 -312 346 -310
rect 366 -312 374 -310
rect 412 -328 414 -306
rect 562 -307 564 -304
rect 379 -334 381 -328
rect 340 -338 342 -335
rect 806 -299 808 -296
rect 412 -371 414 -368
rect 562 -369 564 -347
rect 595 -353 597 -341
rect 671 -358 673 -336
rect 704 -358 706 -336
rect 878 -332 880 -329
rect 839 -339 841 -333
rect 602 -364 610 -362
rect 630 -364 633 -362
rect 379 -377 381 -374
rect 340 -381 342 -378
rect 806 -361 808 -339
rect 846 -357 854 -355
rect 874 -357 877 -355
rect 671 -381 673 -378
rect 704 -381 706 -378
rect 891 -362 893 -358
rect 806 -384 808 -381
rect 891 -385 893 -382
rect 562 -392 564 -389
<< polycontact >>
rect 245 666 249 670
rect 685 647 689 651
rect 718 647 722 651
rect 751 647 755 651
rect 784 647 788 651
rect 817 647 821 651
rect 852 646 856 650
rect 515 618 519 622
rect 548 618 552 622
rect 581 618 585 622
rect 614 618 618 622
rect 649 617 653 621
rect 200 580 204 584
rect 236 588 240 592
rect 309 591 313 595
rect 342 591 346 595
rect 378 597 382 601
rect 411 597 415 601
rect 444 597 448 601
rect 479 596 483 600
rect 788 619 794 625
rect 240 580 244 584
rect 415 569 421 575
rect 585 590 591 596
rect 788 600 794 606
rect 788 581 794 587
rect 585 571 591 577
rect 788 562 794 568
rect 415 550 421 556
rect 585 552 591 558
rect 788 543 794 549
rect 257 528 261 532
rect 415 531 421 537
rect 585 533 591 539
rect 878 528 882 532
rect 725 523 729 527
rect 877 495 881 499
rect 724 489 728 493
rect 212 442 216 446
rect 248 450 252 454
rect 321 453 325 457
rect 354 453 358 457
rect 394 455 398 459
rect 427 455 431 459
rect 460 455 464 459
rect 495 454 499 458
rect 531 457 535 461
rect 564 457 568 461
rect 597 457 601 461
rect 630 457 634 461
rect 665 456 669 460
rect 876 461 880 465
rect 724 454 728 458
rect 252 442 256 446
rect 431 427 437 433
rect 601 429 607 435
rect 431 408 437 414
rect 601 410 607 416
rect 876 426 880 430
rect 774 414 778 418
rect 690 401 694 405
rect 711 401 715 405
rect 740 401 744 405
rect 774 401 778 405
rect 797 402 801 406
rect 310 390 314 394
rect 431 389 437 395
rect 601 391 607 397
rect 601 373 607 379
rect 926 386 930 390
rect 822 373 826 377
rect 842 373 846 377
rect 863 373 867 377
rect 892 373 896 377
rect 926 373 930 377
rect 949 374 953 378
rect 265 304 269 308
rect 301 312 305 316
rect 374 315 378 319
rect 407 315 411 319
rect 610 350 614 354
rect 768 325 772 329
rect 610 315 614 319
rect 305 304 309 308
rect 450 294 454 298
rect 483 294 487 298
rect 516 294 520 298
rect 551 293 555 297
rect 487 266 493 272
rect 660 275 664 279
rect 597 262 601 266
rect 626 262 630 266
rect 660 262 664 266
rect 683 263 687 267
rect 806 278 812 283
rect 310 252 314 256
rect 487 247 493 253
rect 732 258 736 262
rect 841 269 845 273
rect 874 269 878 273
rect 772 257 776 261
rect 819 257 825 262
rect 487 228 493 234
rect 265 166 269 170
rect 301 174 305 178
rect 374 177 378 181
rect 407 177 411 181
rect 438 177 442 181
rect 305 166 309 170
rect 488 137 492 141
rect 454 124 458 128
rect 488 124 492 128
rect 511 125 515 129
rect 603 135 607 139
rect 324 88 330 93
rect 373 89 377 93
rect 271 77 275 81
rect 304 77 308 81
rect 413 88 417 92
rect 337 67 343 72
rect 558 49 562 53
rect 594 57 598 61
rect 667 60 671 64
rect 700 60 704 64
rect 598 49 602 53
rect 377 21 381 25
rect 600 -3 604 1
rect 324 -46 330 -41
rect 373 -45 377 -41
rect 271 -57 275 -53
rect 304 -57 308 -53
rect 413 -46 417 -42
rect 337 -67 343 -62
rect 828 -22 832 -18
rect 555 -89 559 -85
rect 591 -81 595 -77
rect 664 -78 668 -74
rect 697 -78 701 -74
rect 866 -69 872 -64
rect 595 -89 599 -85
rect 377 -113 381 -109
rect 792 -89 796 -85
rect 832 -90 836 -86
rect 879 -90 885 -85
rect 603 -141 607 -137
rect 825 -156 829 -152
rect 325 -180 331 -175
rect 374 -179 378 -175
rect 414 -180 418 -176
rect 338 -201 344 -196
rect 558 -227 562 -223
rect 863 -203 869 -198
rect 594 -219 598 -215
rect 789 -223 793 -219
rect 598 -227 602 -223
rect 829 -224 833 -220
rect 876 -224 882 -219
rect 378 -247 382 -243
rect 603 -279 607 -275
rect 838 -290 842 -286
rect 325 -314 331 -309
rect 374 -313 378 -309
rect 414 -314 418 -310
rect 338 -335 344 -330
rect 558 -365 562 -361
rect 594 -357 598 -353
rect 667 -354 671 -350
rect 700 -354 704 -350
rect 876 -337 882 -332
rect 802 -357 806 -353
rect 598 -365 602 -361
rect 378 -381 382 -377
rect 842 -358 846 -354
rect 889 -358 895 -353
<< metal1 >>
rect 663 714 869 717
rect 663 713 699 714
rect 663 688 666 713
rect 675 710 699 713
rect 708 710 732 714
rect 741 710 765 714
rect 774 710 798 714
rect 807 710 831 714
rect 845 710 869 714
rect 493 685 666 688
rect 493 684 529 685
rect 272 670 285 674
rect 185 666 245 670
rect 185 584 190 666
rect 268 653 272 662
rect 193 644 217 651
rect 226 650 272 653
rect 232 644 236 650
rect 199 638 203 644
rect 207 584 211 598
rect 240 599 244 604
rect 279 599 285 670
rect 493 667 496 684
rect 505 681 529 684
rect 538 681 562 685
rect 571 681 595 685
rect 604 681 628 685
rect 642 681 666 685
rect 681 704 685 710
rect 714 704 718 710
rect 747 704 751 710
rect 780 704 784 710
rect 813 704 817 710
rect 851 704 855 710
rect 356 664 496 667
rect 356 663 392 664
rect 356 662 359 663
rect 302 655 359 662
rect 368 660 392 663
rect 401 660 425 664
rect 434 660 458 664
rect 472 660 496 664
rect 511 675 515 681
rect 544 675 548 681
rect 577 675 581 681
rect 610 675 614 681
rect 648 675 652 681
rect 308 649 312 655
rect 341 649 345 655
rect 374 654 378 660
rect 407 654 411 660
rect 440 654 444 660
rect 478 654 482 660
rect 689 654 693 664
rect 722 654 726 664
rect 755 654 759 664
rect 788 654 792 664
rect 821 654 825 664
rect 519 625 523 635
rect 552 625 556 635
rect 585 625 589 635
rect 618 625 622 635
rect 240 596 285 599
rect 240 595 302 596
rect 316 595 320 609
rect 349 595 353 609
rect 382 604 386 614
rect 415 604 419 614
rect 448 604 452 614
rect 236 584 240 588
rect 272 584 276 595
rect 282 591 309 595
rect 316 591 342 595
rect 349 591 361 595
rect 316 587 320 591
rect 349 587 353 591
rect 185 580 200 584
rect 207 580 240 584
rect 185 -321 188 580
rect 207 576 211 580
rect 199 547 203 556
rect 268 547 272 576
rect 308 547 312 567
rect 341 547 345 567
rect 193 539 360 547
rect 378 537 382 597
rect 401 597 411 601
rect 486 600 490 614
rect 401 556 405 597
rect 444 592 448 597
rect 415 589 448 592
rect 460 596 479 600
rect 486 596 501 600
rect 415 575 421 589
rect 460 578 464 596
rect 486 592 490 596
rect 478 570 482 572
rect 460 559 464 566
rect 401 550 415 556
rect 472 567 482 570
rect 460 540 464 547
rect 284 532 297 536
rect 196 528 257 532
rect 196 446 202 528
rect 280 515 284 524
rect 205 506 229 513
rect 238 512 284 515
rect 244 506 248 512
rect 277 511 284 512
rect 211 500 215 506
rect 219 446 223 460
rect 252 461 256 466
rect 291 461 297 532
rect 378 531 415 537
rect 472 532 476 567
rect 515 539 519 618
rect 548 558 552 618
rect 571 618 581 622
rect 656 621 660 635
rect 571 577 575 618
rect 614 613 618 618
rect 585 610 618 613
rect 630 617 649 621
rect 656 617 671 621
rect 585 596 591 610
rect 630 599 634 617
rect 656 613 660 617
rect 648 591 652 593
rect 630 580 634 587
rect 571 571 585 577
rect 642 588 652 591
rect 630 561 634 568
rect 548 552 585 558
rect 630 542 634 549
rect 515 533 585 539
rect 642 534 646 588
rect 685 549 689 647
rect 718 568 722 647
rect 751 587 755 647
rect 774 647 784 651
rect 859 650 863 664
rect 774 606 778 647
rect 817 642 821 647
rect 788 639 821 642
rect 833 646 852 650
rect 859 646 874 650
rect 788 625 794 639
rect 833 628 837 646
rect 859 642 863 646
rect 851 620 855 622
rect 833 609 837 616
rect 774 600 788 606
rect 845 617 855 620
rect 833 590 837 597
rect 751 581 788 587
rect 833 571 837 578
rect 718 562 788 568
rect 833 552 837 559
rect 685 543 788 549
rect 845 544 849 617
rect 837 540 849 544
rect 464 528 476 532
rect 634 530 646 534
rect 925 532 947 536
rect 772 527 795 531
rect 521 525 682 527
rect 384 524 682 525
rect 314 522 545 524
rect 314 521 408 522
rect 314 517 371 521
rect 384 518 408 521
rect 417 518 441 522
rect 450 518 474 522
rect 488 518 512 522
rect 521 520 545 522
rect 554 520 578 524
rect 587 520 611 524
rect 620 520 644 524
rect 658 520 682 524
rect 690 523 725 527
rect 320 511 324 517
rect 353 511 357 517
rect 390 512 394 518
rect 423 512 427 518
rect 456 512 460 518
rect 494 512 498 518
rect 527 514 531 520
rect 560 514 564 520
rect 593 514 597 520
rect 626 514 630 520
rect 664 514 668 520
rect 252 458 297 461
rect 252 457 314 458
rect 328 457 332 471
rect 361 457 365 471
rect 398 462 402 472
rect 431 462 435 472
rect 464 462 468 472
rect 248 446 252 450
rect 284 446 288 457
rect 294 453 321 457
rect 328 453 354 457
rect 361 453 373 457
rect 328 449 332 453
rect 361 449 365 453
rect 196 442 212 446
rect 219 442 252 446
rect 196 -186 203 442
rect 219 438 223 442
rect 211 409 215 418
rect 280 409 284 438
rect 320 409 324 429
rect 353 409 357 429
rect 208 401 372 409
rect 337 394 350 398
rect 250 390 310 394
rect 250 308 255 390
rect 333 377 337 386
rect 258 368 282 375
rect 291 374 337 377
rect 297 368 301 374
rect 264 362 268 368
rect 272 308 276 322
rect 305 323 309 328
rect 344 323 350 394
rect 394 395 398 455
rect 417 455 427 459
rect 502 458 506 472
rect 535 464 539 474
rect 568 464 572 474
rect 601 464 605 474
rect 634 464 638 474
rect 417 414 421 455
rect 460 450 464 455
rect 431 447 464 450
rect 476 454 495 458
rect 502 454 517 458
rect 431 433 437 447
rect 476 436 480 454
rect 502 450 506 454
rect 494 428 498 430
rect 476 417 480 424
rect 417 408 431 414
rect 488 425 498 428
rect 476 398 480 405
rect 394 389 431 395
rect 488 390 492 425
rect 480 386 492 390
rect 367 379 424 386
rect 531 379 535 457
rect 564 397 568 457
rect 587 457 597 461
rect 672 460 676 474
rect 587 416 591 457
rect 630 452 634 457
rect 601 449 634 452
rect 646 456 665 460
rect 672 456 687 460
rect 601 435 607 449
rect 646 438 650 456
rect 672 452 676 456
rect 664 430 668 432
rect 646 419 650 426
rect 587 410 601 416
rect 658 427 668 430
rect 646 400 650 407
rect 564 391 601 397
rect 646 382 650 388
rect 373 373 377 379
rect 406 373 410 379
rect 531 373 601 379
rect 658 374 662 427
rect 690 405 694 523
rect 767 497 772 519
rect 771 493 772 497
rect 711 489 724 493
rect 711 405 715 489
rect 766 462 771 485
rect 790 473 795 527
rect 822 528 878 532
rect 790 466 814 473
rect 796 460 800 466
rect 720 454 724 458
rect 731 444 735 450
rect 723 440 735 444
rect 723 421 727 440
rect 771 425 787 429
rect 723 417 731 421
rect 740 405 744 409
rect 774 405 778 414
rect 782 406 787 425
rect 804 406 808 420
rect 782 402 797 406
rect 804 402 819 406
rect 698 394 699 398
rect 719 394 720 398
rect 748 394 749 398
rect 781 394 782 398
rect 787 394 791 402
rect 804 398 808 402
rect 686 374 690 378
rect 707 374 711 378
rect 736 374 740 378
rect 769 374 773 378
rect 796 374 800 378
rect 650 371 800 374
rect 822 377 826 528
rect 920 503 925 524
rect 924 499 925 503
rect 842 495 877 499
rect 842 377 846 495
rect 919 469 924 491
rect 923 465 924 469
rect 863 461 876 465
rect 863 377 867 461
rect 918 434 923 457
rect 942 445 947 532
rect 942 438 966 445
rect 948 432 952 438
rect 872 426 876 430
rect 883 416 887 422
rect 875 412 887 416
rect 875 393 879 412
rect 923 397 939 401
rect 875 389 883 393
rect 892 377 896 379
rect 926 377 930 386
rect 934 378 939 397
rect 956 378 960 392
rect 934 374 949 378
rect 956 374 971 378
rect 650 370 662 371
rect 440 361 568 364
rect 440 357 464 361
rect 473 357 497 361
rect 506 357 530 361
rect 544 357 568 361
rect 305 320 350 323
rect 305 319 367 320
rect 381 319 385 333
rect 414 319 418 333
rect 446 351 450 357
rect 479 351 483 357
rect 512 351 516 357
rect 550 351 554 357
rect 657 354 681 358
rect 301 308 305 312
rect 337 308 341 319
rect 347 315 374 319
rect 381 315 407 319
rect 414 315 426 319
rect 381 311 385 315
rect 414 311 418 315
rect 209 304 265 308
rect 272 304 305 308
rect 209 -53 216 304
rect 272 300 276 304
rect 264 271 268 280
rect 333 271 337 300
rect 454 301 458 311
rect 487 301 491 311
rect 520 301 524 311
rect 373 271 377 291
rect 406 271 410 291
rect 257 263 424 271
rect 337 256 350 260
rect 250 252 310 256
rect 250 170 255 252
rect 333 239 337 248
rect 258 230 282 237
rect 291 236 337 239
rect 297 230 301 236
rect 264 224 268 230
rect 272 170 276 184
rect 305 185 309 190
rect 344 185 350 256
rect 367 241 424 248
rect 373 235 377 241
rect 406 235 410 241
rect 450 234 454 294
rect 473 294 483 298
rect 558 297 562 311
rect 597 350 610 354
rect 473 253 477 294
rect 516 289 520 294
rect 487 286 520 289
rect 532 293 551 297
rect 558 293 573 297
rect 487 272 493 286
rect 532 275 536 293
rect 558 289 562 293
rect 550 267 554 269
rect 532 256 536 263
rect 473 247 487 253
rect 544 264 554 267
rect 597 266 601 350
rect 652 323 657 346
rect 676 334 681 354
rect 830 366 831 370
rect 850 366 851 370
rect 871 366 872 370
rect 900 366 901 370
rect 933 366 934 370
rect 939 366 943 374
rect 956 370 960 374
rect 717 344 807 348
rect 676 327 700 334
rect 682 321 686 327
rect 607 315 610 319
rect 617 305 621 311
rect 609 301 621 305
rect 609 282 613 301
rect 657 286 673 290
rect 609 278 617 282
rect 532 237 536 244
rect 450 228 487 234
rect 544 229 548 264
rect 626 266 630 269
rect 660 266 664 275
rect 668 267 673 286
rect 690 267 694 281
rect 668 263 683 267
rect 690 263 705 267
rect 605 255 606 259
rect 634 255 635 259
rect 667 255 668 259
rect 673 255 677 263
rect 690 259 694 263
rect 717 262 722 344
rect 768 329 772 344
rect 725 322 749 329
rect 803 326 807 344
rect 818 346 822 350
rect 838 346 842 350
rect 859 346 863 350
rect 888 346 892 350
rect 921 346 925 350
rect 948 346 952 350
rect 818 343 952 346
rect 834 333 891 340
rect 840 327 844 333
rect 873 327 877 333
rect 731 316 735 322
rect 739 262 743 276
rect 717 258 732 262
rect 739 258 754 262
rect 739 254 743 258
rect 593 235 597 239
rect 622 235 626 239
rect 655 235 659 239
rect 682 235 686 239
rect 593 232 686 235
rect 749 248 754 258
rect 764 261 768 282
rect 815 286 833 290
rect 772 273 776 282
rect 806 276 812 278
rect 829 273 833 286
rect 848 273 852 287
rect 881 273 885 287
rect 772 269 841 273
rect 848 269 874 273
rect 881 269 893 273
rect 804 261 807 269
rect 764 257 772 261
rect 810 258 819 261
rect 784 248 788 253
rect 810 248 813 258
rect 749 245 813 248
rect 749 244 788 245
rect 536 225 548 229
rect 731 225 735 234
rect 831 250 835 269
rect 848 265 852 269
rect 881 265 885 269
rect 828 247 835 250
rect 840 225 844 245
rect 873 225 877 245
rect 725 217 892 225
rect 305 182 350 185
rect 305 181 367 182
rect 381 181 385 195
rect 414 181 418 195
rect 480 191 528 196
rect 480 185 485 191
rect 504 189 528 191
rect 510 183 514 189
rect 301 170 305 174
rect 337 170 341 181
rect 347 177 374 181
rect 381 177 407 181
rect 414 177 438 181
rect 381 173 385 177
rect 414 173 418 177
rect 238 166 265 170
rect 272 166 305 170
rect 238 81 243 166
rect 272 162 276 166
rect 264 133 268 142
rect 333 133 337 162
rect 373 133 377 153
rect 406 133 410 153
rect 257 125 424 133
rect 427 128 431 177
rect 445 167 449 173
rect 437 163 449 167
rect 437 144 441 163
rect 485 148 501 152
rect 437 140 445 144
rect 488 128 492 137
rect 272 105 276 125
rect 305 105 309 125
rect 314 100 321 103
rect 264 81 268 85
rect 297 81 301 85
rect 314 81 318 100
rect 414 116 418 125
rect 427 124 454 128
rect 496 129 501 148
rect 518 129 522 143
rect 630 139 643 143
rect 543 135 603 139
rect 496 125 511 129
rect 518 125 533 129
rect 361 105 400 106
rect 336 102 400 105
rect 336 92 339 102
rect 361 97 365 102
rect 330 89 339 92
rect 377 89 385 93
rect 342 81 345 89
rect 238 77 268 81
rect 275 77 301 81
rect 308 77 377 81
rect 264 63 268 77
rect 297 63 301 77
rect 316 64 320 77
rect 337 72 343 74
rect 373 68 377 77
rect 316 60 334 64
rect 381 68 385 89
rect 395 92 400 102
rect 462 117 463 121
rect 495 117 496 121
rect 501 117 505 125
rect 518 121 522 125
rect 450 97 454 101
rect 483 97 487 101
rect 510 97 514 101
rect 406 92 410 96
rect 448 94 514 97
rect 395 88 410 92
rect 417 88 432 92
rect 406 74 410 88
rect 414 28 418 34
rect 427 38 432 88
rect 543 53 548 135
rect 626 122 630 131
rect 551 113 575 120
rect 584 119 630 122
rect 590 113 594 119
rect 557 107 561 113
rect 565 53 569 67
rect 598 68 602 73
rect 637 68 643 139
rect 660 124 717 131
rect 666 118 670 124
rect 699 118 703 124
rect 598 65 643 68
rect 598 64 660 65
rect 674 64 678 78
rect 707 64 711 78
rect 594 53 598 57
rect 630 53 634 64
rect 640 60 667 64
rect 674 60 700 64
rect 707 60 719 64
rect 674 56 678 60
rect 707 56 711 60
rect 743 58 762 66
rect 543 49 558 53
rect 565 49 598 53
rect 565 45 569 49
rect 427 30 505 38
rect 272 17 276 23
rect 305 17 309 23
rect 258 10 315 17
rect 342 6 346 24
rect 400 21 424 28
rect 377 6 381 21
rect 427 6 432 30
rect 470 25 505 30
rect 470 9 505 22
rect 557 16 561 25
rect 626 16 630 45
rect 666 16 670 36
rect 699 16 703 36
rect 551 8 718 16
rect 342 2 432 6
rect 627 1 640 5
rect 257 -9 424 -1
rect 540 -3 600 1
rect 272 -29 276 -9
rect 305 -29 309 -9
rect 314 -34 321 -31
rect 264 -53 268 -49
rect 297 -53 301 -49
rect 314 -53 318 -34
rect 414 -18 418 -9
rect 361 -29 400 -28
rect 336 -32 400 -29
rect 336 -42 339 -32
rect 361 -37 365 -32
rect 330 -45 339 -42
rect 377 -45 385 -41
rect 342 -53 345 -45
rect 209 -57 268 -53
rect 275 -57 301 -53
rect 308 -57 377 -53
rect 264 -71 268 -57
rect 297 -71 301 -57
rect 316 -70 320 -57
rect 337 -62 343 -60
rect 373 -66 377 -57
rect 316 -74 334 -70
rect 381 -66 385 -45
rect 395 -42 400 -32
rect 406 -42 410 -38
rect 395 -46 410 -42
rect 417 -46 432 -42
rect 406 -60 410 -46
rect 414 -106 418 -100
rect 427 -101 432 -46
rect 540 -85 545 -3
rect 623 -16 627 -7
rect 548 -25 572 -18
rect 581 -19 627 -16
rect 587 -25 591 -19
rect 554 -31 558 -25
rect 562 -85 566 -71
rect 595 -70 599 -65
rect 634 -70 640 1
rect 777 -3 867 1
rect 657 -14 714 -7
rect 663 -20 667 -14
rect 696 -20 700 -14
rect 595 -73 640 -70
rect 595 -74 657 -73
rect 671 -74 675 -60
rect 704 -74 708 -60
rect 591 -85 595 -81
rect 627 -85 631 -74
rect 637 -78 664 -74
rect 671 -78 697 -74
rect 704 -78 716 -74
rect 671 -82 675 -78
rect 704 -82 708 -78
rect 744 -80 756 -72
rect 540 -89 555 -85
rect 562 -89 595 -85
rect 562 -93 566 -89
rect 470 -101 505 -99
rect 272 -117 276 -111
rect 305 -117 309 -111
rect 258 -124 315 -117
rect 342 -128 346 -110
rect 400 -113 424 -106
rect 427 -107 505 -101
rect 377 -128 381 -113
rect 427 -128 432 -107
rect 470 -112 505 -107
rect 470 -127 505 -115
rect 554 -122 558 -113
rect 623 -122 627 -93
rect 777 -85 782 -3
rect 828 -18 832 -3
rect 785 -25 809 -18
rect 863 -21 867 -3
rect 791 -31 795 -25
rect 799 -85 803 -71
rect 777 -89 792 -85
rect 799 -89 814 -85
rect 799 -93 803 -89
rect 663 -122 667 -102
rect 696 -122 700 -102
rect 809 -99 814 -89
rect 824 -86 828 -65
rect 875 -61 893 -57
rect 832 -74 836 -65
rect 866 -71 872 -69
rect 889 -74 893 -61
rect 832 -78 894 -74
rect 864 -86 867 -78
rect 824 -90 832 -86
rect 870 -89 879 -86
rect 844 -99 848 -94
rect 870 -99 873 -89
rect 809 -102 873 -99
rect 809 -103 848 -102
rect 791 -122 795 -113
rect 891 -97 894 -78
rect 888 -100 894 -97
rect 342 -132 432 -128
rect 548 -130 715 -122
rect 785 -130 894 -122
rect 317 -143 425 -135
rect 630 -137 643 -133
rect 543 -141 603 -137
rect 315 -168 322 -165
rect 315 -186 319 -168
rect 415 -152 419 -143
rect 362 -163 401 -162
rect 337 -166 401 -163
rect 337 -176 340 -166
rect 362 -171 366 -166
rect 331 -179 340 -176
rect 378 -179 386 -175
rect 196 -187 319 -186
rect 343 -187 346 -179
rect 196 -191 378 -187
rect 317 -204 321 -191
rect 338 -196 344 -194
rect 374 -200 378 -191
rect 317 -208 335 -204
rect 382 -200 386 -179
rect 396 -176 401 -166
rect 407 -176 411 -172
rect 396 -180 411 -176
rect 418 -180 433 -176
rect 407 -194 411 -180
rect 415 -240 419 -234
rect 428 -240 433 -180
rect 543 -223 548 -141
rect 626 -154 630 -145
rect 551 -163 575 -156
rect 584 -157 630 -154
rect 590 -163 594 -157
rect 557 -169 561 -163
rect 565 -223 569 -209
rect 598 -208 602 -203
rect 637 -208 643 -137
rect 598 -211 643 -208
rect 774 -137 864 -133
rect 774 -211 779 -137
rect 825 -152 829 -137
rect 782 -159 806 -152
rect 860 -155 864 -137
rect 788 -165 792 -159
rect 598 -212 766 -211
rect 594 -223 598 -219
rect 630 -223 634 -212
rect 640 -216 766 -212
rect 660 -217 766 -216
rect 746 -219 766 -217
rect 771 -219 779 -211
rect 796 -219 800 -205
rect 774 -223 789 -219
rect 796 -223 811 -219
rect 543 -227 558 -223
rect 565 -227 598 -223
rect 796 -227 800 -223
rect 565 -231 569 -227
rect 470 -240 505 -237
rect 343 -262 347 -244
rect 401 -247 425 -240
rect 428 -246 505 -240
rect 378 -262 382 -247
rect 428 -262 433 -246
rect 470 -249 505 -246
rect 343 -266 433 -262
rect 470 -265 505 -252
rect 557 -260 561 -251
rect 626 -260 630 -231
rect 806 -233 811 -223
rect 821 -220 825 -199
rect 872 -195 890 -191
rect 829 -208 833 -199
rect 863 -205 869 -203
rect 886 -208 890 -195
rect 829 -212 891 -208
rect 861 -220 864 -212
rect 821 -224 829 -220
rect 867 -223 876 -220
rect 841 -233 845 -228
rect 867 -233 870 -223
rect 806 -236 870 -233
rect 806 -237 845 -236
rect 788 -256 792 -247
rect 888 -231 891 -212
rect 885 -234 891 -231
rect 551 -268 660 -260
rect 782 -264 891 -256
rect 317 -277 425 -269
rect 787 -271 877 -267
rect 630 -275 643 -271
rect 315 -302 322 -299
rect 315 -321 319 -302
rect 415 -286 419 -277
rect 362 -297 401 -296
rect 337 -300 401 -297
rect 337 -310 340 -300
rect 362 -305 366 -300
rect 331 -313 340 -310
rect 378 -313 386 -309
rect 343 -321 346 -313
rect 185 -325 378 -321
rect 256 -326 322 -325
rect 317 -338 321 -326
rect 338 -330 344 -328
rect 374 -334 378 -325
rect 317 -342 335 -338
rect 317 -425 320 -342
rect 382 -334 386 -313
rect 396 -310 401 -300
rect 543 -279 603 -275
rect 407 -310 411 -306
rect 396 -314 411 -310
rect 418 -314 433 -310
rect 407 -328 411 -314
rect 415 -374 419 -368
rect 343 -396 347 -378
rect 401 -381 425 -374
rect 378 -396 382 -381
rect 428 -382 433 -314
rect 543 -361 548 -279
rect 626 -292 630 -283
rect 551 -301 575 -294
rect 584 -295 630 -292
rect 590 -301 594 -295
rect 557 -307 561 -301
rect 565 -361 569 -347
rect 598 -346 602 -341
rect 637 -346 643 -275
rect 660 -290 717 -283
rect 666 -296 670 -290
rect 699 -296 703 -290
rect 598 -349 643 -346
rect 598 -350 660 -349
rect 674 -350 678 -336
rect 707 -350 711 -336
rect 594 -361 598 -357
rect 630 -361 634 -350
rect 640 -354 667 -350
rect 674 -354 700 -350
rect 707 -354 719 -350
rect 674 -358 678 -354
rect 707 -358 711 -354
rect 746 -356 774 -348
rect 787 -353 792 -271
rect 838 -286 842 -271
rect 795 -293 819 -286
rect 873 -289 877 -271
rect 801 -299 805 -293
rect 809 -353 813 -339
rect 543 -365 558 -361
rect 565 -365 598 -361
rect 565 -369 569 -365
rect 470 -382 505 -377
rect 428 -388 505 -382
rect 428 -396 433 -388
rect 470 -390 505 -388
rect 343 -400 433 -396
rect 470 -406 505 -393
rect 557 -398 561 -389
rect 626 -398 630 -369
rect 787 -357 802 -353
rect 809 -357 824 -353
rect 666 -398 670 -378
rect 699 -398 703 -378
rect 551 -406 718 -398
rect 787 -404 791 -357
rect 809 -361 813 -357
rect 819 -367 824 -357
rect 834 -354 838 -333
rect 885 -329 903 -325
rect 842 -342 846 -333
rect 876 -339 882 -337
rect 899 -342 903 -329
rect 842 -346 905 -342
rect 874 -354 877 -346
rect 834 -358 842 -354
rect 880 -357 889 -354
rect 854 -367 858 -362
rect 880 -367 883 -357
rect 819 -370 883 -367
rect 819 -371 858 -370
rect 801 -390 805 -381
rect 901 -365 905 -346
rect 898 -368 905 -365
rect 795 -398 905 -390
rect 787 -414 794 -404
rect 790 -425 794 -414
rect 317 -428 794 -425
<< metal2 >>
rect 208 655 302 662
rect 208 651 216 655
rect 694 654 722 659
rect 727 654 755 659
rect 760 654 788 659
rect 793 654 821 659
rect 826 654 842 659
rect 838 651 842 654
rect 265 607 272 644
rect 524 625 552 630
rect 557 625 585 630
rect 590 625 618 630
rect 623 625 639 630
rect 635 622 639 625
rect 172 603 272 607
rect 387 604 415 609
rect 420 604 448 609
rect 453 604 469 609
rect 172 -267 177 603
rect 465 601 469 604
rect 220 517 314 524
rect 220 513 228 517
rect 277 483 284 505
rect 181 477 284 483
rect 181 -128 192 477
rect 403 462 431 467
rect 436 462 464 467
rect 469 462 485 467
rect 540 464 568 469
rect 573 464 601 469
rect 606 464 634 469
rect 639 464 655 469
rect 481 459 485 462
rect 651 461 655 464
rect 715 409 719 458
rect 715 405 740 409
rect 699 394 715 398
rect 720 394 744 398
rect 749 394 777 398
rect 782 394 787 398
rect 273 379 367 386
rect 867 381 871 430
rect 273 375 281 379
rect 867 377 892 381
rect 337 368 576 373
rect 459 301 487 306
rect 492 301 520 306
rect 525 301 541 306
rect 537 298 541 301
rect 273 241 367 248
rect 273 237 281 241
rect 572 165 576 368
rect 831 366 846 370
rect 851 366 867 370
rect 872 366 896 370
rect 901 366 929 370
rect 934 366 939 370
rect 740 333 834 340
rect 740 329 748 333
rect 601 270 605 319
rect 806 271 812 276
rect 601 266 626 270
rect 769 265 812 271
rect 606 255 630 259
rect 635 255 663 259
rect 668 255 673 259
rect 807 232 812 265
rect 488 160 733 165
rect 488 135 492 160
rect 566 126 660 131
rect 337 85 342 118
rect 463 117 491 121
rect 496 117 501 121
rect 566 120 574 126
rect 337 79 381 85
rect 386 79 463 85
rect 337 73 343 79
rect 455 21 463 79
rect 615 21 620 114
rect 727 66 733 160
rect 720 58 740 66
rect 401 17 409 21
rect 315 10 409 17
rect 455 14 494 21
rect 502 16 620 21
rect 563 -12 657 -7
rect 337 -49 342 -16
rect 563 -18 571 -12
rect 337 -55 381 -49
rect 386 -55 452 -49
rect 337 -60 343 -55
rect 401 -117 409 -113
rect 315 -124 409 -117
rect 443 -116 452 -55
rect 610 -116 617 -23
rect 720 -80 741 -72
rect 866 -76 872 -71
rect 443 -123 491 -116
rect 501 -121 617 -116
rect 728 -128 735 -80
rect 829 -82 872 -76
rect 867 -115 872 -82
rect 181 -135 735 -128
rect 338 -183 343 -150
rect 338 -189 382 -183
rect 387 -189 451 -183
rect 338 -194 344 -189
rect 444 -254 451 -189
rect 619 -254 624 -161
rect 863 -210 869 -205
rect 723 -219 743 -211
rect 826 -216 869 -210
rect 444 -259 496 -254
rect 503 -259 624 -254
rect 731 -267 739 -219
rect 864 -249 869 -216
rect 172 -268 660 -267
rect 719 -268 739 -267
rect 172 -272 739 -268
rect 338 -317 343 -284
rect 566 -287 660 -283
rect 566 -294 574 -287
rect 338 -323 382 -317
rect 387 -323 450 -317
rect 338 -328 344 -323
rect 442 -394 450 -323
rect 617 -393 622 -299
rect 876 -344 882 -339
rect 723 -356 743 -348
rect 839 -350 882 -344
rect 877 -383 882 -350
rect 442 -400 496 -394
rect 503 -397 622 -393
<< metal3 >>
rect 489 47 554 55
rect 489 32 496 47
rect 493 -88 553 -82
rect 493 -102 500 -88
rect 496 -229 556 -223
rect 496 -240 503 -229
rect 494 -367 557 -361
rect 494 -379 501 -367
<< metal4 >>
rect 815 277 822 407
rect 815 271 909 277
rect 901 -105 909 271
rect 880 -112 910 -105
rect 315 -224 321 -204
rect 315 -230 537 -224
rect 531 -239 537 -230
rect 773 -239 779 -218
rect 531 -246 779 -239
rect 881 -274 889 -112
rect 834 -282 889 -274
rect 834 -350 843 -282
<< pad >>
rect 302 655 310 662
rect 689 654 694 659
rect 722 654 727 659
rect 755 654 760 659
rect 788 654 793 659
rect 821 654 826 659
rect 208 644 216 651
rect 265 644 272 651
rect 838 646 843 651
rect 519 625 524 630
rect 552 625 557 630
rect 585 625 590 630
rect 618 625 623 630
rect 635 617 640 622
rect 382 604 387 609
rect 415 604 420 609
rect 448 604 453 609
rect 465 596 470 601
rect 314 517 322 524
rect 220 506 228 513
rect 277 505 284 512
rect 398 462 403 467
rect 431 462 436 467
rect 464 462 469 467
rect 535 464 540 469
rect 568 464 573 469
rect 601 464 606 469
rect 634 464 639 469
rect 481 454 486 459
rect 651 456 656 461
rect 719 454 724 459
rect 871 426 876 431
rect 740 405 745 410
rect 815 402 820 407
rect 694 394 699 399
rect 715 394 720 399
rect 744 394 749 399
rect 777 394 782 399
rect 787 394 792 399
rect 367 379 375 386
rect 892 377 897 382
rect 273 368 281 375
rect 330 368 337 375
rect 826 366 831 371
rect 846 366 851 371
rect 867 366 872 371
rect 896 366 901 371
rect 929 366 934 371
rect 939 366 944 371
rect 834 333 842 340
rect 740 322 748 329
rect 605 315 610 320
rect 454 301 459 306
rect 487 301 492 306
rect 520 301 525 306
rect 537 293 542 298
rect 806 276 812 281
rect 626 266 631 271
rect 764 265 769 271
rect 601 255 606 260
rect 630 255 635 260
rect 663 255 668 260
rect 673 255 678 260
rect 367 241 375 248
rect 273 230 281 237
rect 812 233 818 238
rect 488 130 493 135
rect 660 124 668 131
rect 332 113 337 118
rect 458 117 463 122
rect 491 117 496 122
rect 501 117 506 122
rect 566 113 574 120
rect 615 114 623 122
rect 381 79 386 85
rect 337 70 343 76
rect 712 58 720 66
rect 740 58 748 66
rect 554 47 562 55
rect 489 30 497 38
rect 401 21 409 28
rect 307 10 315 17
rect 494 14 502 22
rect 657 -14 665 -7
rect 332 -21 338 -16
rect 563 -25 571 -18
rect 610 -23 617 -16
rect 800 -25 808 -18
rect 381 -55 386 -49
rect 337 -63 343 -58
rect 866 -71 872 -66
rect 712 -80 720 -72
rect 741 -80 749 -72
rect 824 -82 829 -76
rect 552 -90 559 -83
rect 401 -113 409 -106
rect 491 -108 501 -99
rect 871 -114 877 -109
rect 307 -124 315 -117
rect 491 -124 501 -115
rect 333 -155 339 -150
rect 566 -163 574 -156
rect 619 -161 626 -154
rect 797 -159 805 -152
rect 382 -189 387 -183
rect 338 -197 344 -192
rect 315 -209 321 -204
rect 863 -205 869 -200
rect 719 -218 724 -211
rect 743 -219 751 -211
rect 821 -216 826 -210
rect 555 -229 562 -222
rect 773 -224 779 -218
rect 495 -244 502 -237
rect 869 -248 874 -243
rect 496 -259 503 -252
rect 333 -289 339 -284
rect 660 -290 668 -283
rect 566 -301 574 -294
rect 617 -299 624 -292
rect 810 -293 818 -286
rect 382 -323 387 -317
rect 338 -331 344 -326
rect 876 -339 882 -334
rect 716 -356 723 -349
rect 743 -356 751 -348
rect 834 -350 839 -344
rect 555 -367 562 -360
rect 494 -384 501 -377
rect 882 -382 888 -377
rect 496 -400 503 -393
<< labels >>
rlabel metal1 484 32 484 32 1 a0
rlabel metal1 485 15 485 15 1 b0
rlabel metal1 492 -103 492 -103 1 a1
rlabel metal1 493 -243 493 -243 1 a2
rlabel metal1 493 -399 493 -399 1 b3
rlabel metal1 488 -121 488 -121 1 b1
rlabel metal1 418 129 418 129 5 gnd
rlabel metal1 304 15 304 15 1 vdd
rlabel metal1 413 26 413 26 1 vdd
rlabel metal1 261 79 261 79 3 p0
rlabel metal1 261 -55 261 -55 1 p1
rlabel metal1 413 -108 413 -108 1 vdd
rlabel metal1 304 -119 304 -119 1 vdd
rlabel metal1 418 -5 418 -5 5 gnd
rlabel metal1 419 -139 419 -139 5 gnd
rlabel metal1 414 -242 414 -242 1 vdd
rlabel metal1 419 -273 419 -273 5 gnd
rlabel metal1 414 -376 414 -376 1 vdd
rlabel metal1 411 243 411 243 5 vdd
rlabel metal1 378 243 378 243 5 vdd
rlabel metal1 269 232 269 232 5 vdd
rlabel metal1 332 237 332 237 1 cin
rlabel metal1 422 178 422 178 1 pocin
rlabel metal1 517 193 517 193 5 vdd
rlabel metal1 511 98 511 98 1 gnd
rlabel metal1 530 127 530 127 1 c1
rlabel metal1 418 267 418 267 5 gnd
rlabel metal1 411 381 411 381 5 vdd
rlabel metal1 378 381 378 381 5 vdd
rlabel metal1 269 370 269 370 5 vdd
rlabel metal1 424 317 424 317 1 p1g0
rlabel metal1 545 227 545 227 1 gnd
rlabel metal1 507 363 507 363 5 vdd
rlabel metal1 451 292 451 292 1 p1
rlabel metal1 475 292 475 292 1 p0
rlabel metal1 489 285 489 285 1 cin
rlabel metal1 216 508 216 508 5 vdd
rlabel metal1 358 519 358 519 5 vdd
rlabel metal1 211 405 211 405 1 gnd
rlabel metal1 451 524 451 524 5 vdd
rlabel metal1 489 388 489 388 1 gnd
rlabel metal1 659 390 659 390 1 gnd
rlabel metal1 621 526 621 526 5 vdd
rlabel metal1 797 375 797 375 1 gnd
rlabel metal1 803 470 803 470 5 vdd
rlabel metal1 533 443 533 443 1 p2
rlabel metal1 565 446 565 446 1 p1
rlabel metal1 589 447 589 447 1 p0
rlabel metal1 602 442 602 442 1 cin
rlabel metal1 680 458 680 458 1 p2p1p0c0
rlabel metal1 691 407 691 407 1 g2
rlabel pad 742 408 742 408 1 p2p1p0c0
rlabel metal1 202 444 202 444 3 p2
rlabel metal1 269 514 269 514 1 g1
rlabel metal1 368 454 368 454 1 p2g1
rlabel metal1 396 449 396 449 1 p2
rlabel metal1 418 449 418 449 1 p1
rlabel metal1 434 441 434 441 1 g0
rlabel metal1 511 457 511 457 1 p2p1g0
rlabel metal1 775 409 775 409 1 p2g1
rlabel metal1 204 646 204 646 5 vdd
rlabel metal1 346 657 346 657 5 vdd
rlabel metal1 199 543 199 543 1 gnd
rlabel metal1 435 666 435 666 5 vdd
rlabel metal1 473 530 473 530 1 gnd
rlabel metal1 605 687 605 687 5 vdd
rlabel metal1 643 551 643 551 1 gnd
rlabel metal1 808 716 808 716 5 vdd
rlabel metal1 846 580 846 580 1 gnd
rlabel metal1 949 347 949 347 1 gnd
rlabel metal1 955 442 955 442 5 vdd
rlabel metal1 192 583 192 583 1 p3
rlabel metal1 264 652 264 652 1 g2
rlabel metal1 359 593 359 593 1 p3g2
rlabel metal1 379 591 379 591 1 p3
rlabel metal1 402 591 402 591 1 p2
rlabel metal1 418 585 418 585 1 g1
rlabel metal1 494 597 494 597 1 p3p2g1
rlabel metal1 516 599 516 599 1 p3
rlabel metal1 550 603 550 603 1 p2
rlabel metal1 586 604 586 604 1 g0
rlabel metal1 666 619 666 619 1 p3p2p1g0
rlabel metal1 686 633 686 633 1 p3
rlabel metal1 720 624 720 624 1 p2
rlabel metal1 753 631 753 631 1 p1
rlabel metal1 775 638 775 638 1 p0
rlabel metal1 790 636 790 636 1 cin
rlabel metal1 867 648 867 648 1 p3p2p1p0c0
rlabel metal1 824 398 824 398 1 g3
rlabel metal1 843 395 843 395 1 p3g2
rlabel metal1 864 395 864 395 1 p3p2g1
rlabel metal1 928 379 928 379 1 p3p2p1p0c0
rlabel metal1 966 376 966 376 7 c4
rlabel metal1 736 324 736 324 5 vdd
rlabel metal1 845 335 845 335 5 vdd
rlabel metal1 878 335 878 335 5 vdd
rlabel metal1 731 221 731 221 1 gnd
rlabel metal1 726 260 726 260 1 p0
rlabel pad 766 268 766 268 1 cin
rlabel metal1 892 271 892 271 1 s0
rlabel pad 894 380 894 380 1 p3p2p1g0
rlabel metal1 570 295 570 295 1 p1p0c0
rlabel pad 489 131 489 131 1 g0
rlabel metal1 683 236 683 236 1 gnd
rlabel metal1 689 331 689 331 5 vdd
rlabel metal1 698 265 698 265 1 c2
rlabel metal1 598 272 598 272 1 g1
rlabel pad 628 267 628 267 1 p1g0
rlabel metal1 661 268 661 268 1 p1p0c0
rlabel metal1 573 612 573 612 1 p1
rlabel metal1 712 409 712 409 1 p2p1g0
rlabel metal1 316 -322 316 -322 1 p3
rlabel metal1 319 -189 319 -189 1 p2
rlabel metal1 815 404 815 404 7 c3
rlabel metal1 483 -257 483 -257 1 b2
rlabel metal1 484 -383 484 -383 1 a3
rlabel metal1 562 115 562 115 5 vdd
rlabel metal1 671 126 671 126 5 vdd
rlabel metal1 704 126 704 126 5 vdd
rlabel metal1 619 14 619 14 1 gnd
rlabel metal1 757 62 757 62 1 g0
rlabel metal1 554 -126 554 -126 1 gnd
rlabel metal1 701 -12 701 -12 5 vdd
rlabel metal1 668 -12 668 -12 5 vdd
rlabel metal1 559 -23 559 -23 5 vdd
rlabel metal1 557 -264 557 -264 1 gnd
rlabel metal1 562 -161 562 -161 5 vdd
rlabel metal1 557 -402 557 -402 1 gnd
rlabel metal1 704 -288 704 -288 5 vdd
rlabel metal1 671 -288 671 -288 5 vdd
rlabel metal1 562 -299 562 -299 5 vdd
rlabel metal1 900 -344 900 -344 1 s3
rlabel metal1 836 -343 836 -343 1 c3
rlabel pad 836 -348 836 -348 1 c3
rlabel metal1 791 -356 791 -356 1 p3
rlabel metal1 806 -291 806 -291 5 vdd
rlabel metal1 801 -394 801 -394 1 gnd
rlabel metal1 888 -209 888 -209 1 s2
rlabel pad 823 -213 823 -213 1 c2
rlabel metal1 777 -221 777 -221 1 p2
rlabel metal1 788 -260 788 -260 1 gnd
rlabel metal1 793 -157 793 -157 5 vdd
rlabel metal1 762 -353 762 -353 1 g3
rlabel metal1 761 -212 761 -212 1 g2
rlabel metal1 751 -76 751 -76 1 g1
rlabel metal1 796 -23 796 -23 5 vdd
rlabel metal1 791 -126 791 -126 1 gnd
rlabel metal1 783 -87 783 -87 1 p1
rlabel pad 825 -79 825 -79 1 c1
rlabel metal1 891 -76 891 -76 1 s1
<< end >>
